
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:22:38 03/20/2018 
// Design Name: 
// Module Name:    sine 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sine(Clk,sine_out,cos_out);
    input Clk;
    output [7:0] sine_out,cos_out;
    reg signed [7:0] sine [0:40000];
    reg signed [7:0] cos [0:40000];
  
    integer i;  
    reg [7:0] sine_out,cos_out; 

    initial begin
        i = 0;
cos[0]=78;
cos[1]=78;
cos[2]=78;
cos[3]=78;
cos[4]=78;
cos[5]=78;
cos[6]=78;
cos[7]=78;
cos[8]=78;
cos[9]=78;
cos[10]=78;
cos[11]=78;
cos[12]=78;
cos[13]=78;
cos[14]=78;
cos[15]=78;
cos[16]=78;
cos[17]=78;
cos[18]=78;
cos[19]=78;
cos[20]=78;
cos[21]=78;
cos[22]=78;
cos[23]=78;
cos[24]=78;
cos[25]=78;
cos[26]=78;
cos[27]=78;
cos[28]=78;
cos[29]=78;
cos[30]=78;
cos[31]=78;
cos[32]=78;
cos[33]=78;
cos[34]=78;
cos[35]=78;
cos[36]=78;
cos[37]=78;
cos[38]=78;
cos[39]=78;
cos[40]=78;
cos[41]=78;
cos[42]=78;
cos[43]=78;
cos[44]=78;
cos[45]=78;
cos[46]=78;
cos[47]=78;
cos[48]=78;
cos[49]=78;
cos[50]=78;
cos[51]=78;
cos[52]=78;
cos[53]=78;
cos[54]=78;
cos[55]=78;
cos[56]=78;
cos[57]=78;
cos[58]=78;
cos[59]=78;
cos[60]=78;
cos[61]=78;
cos[62]=78;
cos[63]=78;
cos[64]=78;
cos[65]=78;
cos[66]=78;
cos[67]=78;
cos[68]=78;
cos[69]=78;
cos[70]=78;
cos[71]=78;
cos[72]=78;
cos[73]=78;
cos[74]=78;
cos[75]=78;
cos[76]=78;
cos[77]=78;
cos[78]=78;
cos[79]=78;
cos[80]=78;
cos[81]=78;
cos[82]=78;
cos[83]=78;
cos[84]=78;
cos[85]=78;
cos[86]=78;
cos[87]=78;
cos[88]=78;
cos[89]=78;
cos[90]=78;
cos[91]=78;
cos[92]=78;
cos[93]=78;
cos[94]=78;
cos[95]=78;
cos[96]=78;
cos[97]=78;
cos[98]=78;
cos[99]=78;
cos[100]=78;
cos[101]=78;
cos[102]=78;
cos[103]=78;
cos[104]=78;
cos[105]=78;
cos[106]=78;
cos[107]=78;
cos[108]=78;
cos[109]=78;
cos[110]=78;
cos[111]=78;
cos[112]=78;
cos[113]=78;
cos[114]=78;
cos[115]=78;
cos[116]=78;
cos[117]=78;
cos[118]=78;
cos[119]=78;
cos[120]=78;
cos[121]=78;
cos[122]=78;
cos[123]=78;
cos[124]=78;
cos[125]=78;
cos[126]=78;
cos[127]=78;
cos[128]=78;
cos[129]=78;
cos[130]=78;
cos[131]=78;
cos[132]=78;
cos[133]=78;
cos[134]=78;
cos[135]=78;
cos[136]=78;
cos[137]=78;
cos[138]=78;
cos[139]=78;
cos[140]=78;
cos[141]=78;
cos[142]=78;
cos[143]=78;
cos[144]=78;
cos[145]=78;
cos[146]=78;
cos[147]=78;
cos[148]=78;
cos[149]=78;
cos[150]=78;
cos[151]=78;
cos[152]=78;
cos[153]=78;
cos[154]=78;
cos[155]=78;
cos[156]=78;
cos[157]=78;
cos[158]=78;
cos[159]=78;
cos[160]=78;
cos[161]=78;
cos[162]=78;
cos[163]=78;
cos[164]=78;
cos[165]=78;
cos[166]=78;
cos[167]=78;
cos[168]=78;
cos[169]=78;
cos[170]=78;
cos[171]=78;
cos[172]=78;
cos[173]=78;
cos[174]=78;
cos[175]=78;
cos[176]=78;
cos[177]=78;
cos[178]=78;
cos[179]=78;
cos[180]=78;
cos[181]=78;
cos[182]=78;
cos[183]=78;
cos[184]=78;
cos[185]=78;
cos[186]=78;
cos[187]=78;
cos[188]=78;
cos[189]=78;
cos[190]=78;
cos[191]=78;
cos[192]=78;
cos[193]=78;
cos[194]=78;
cos[195]=78;
cos[196]=78;
cos[197]=78;
cos[198]=78;
cos[199]=78;
cos[200]=78;
cos[201]=78;
cos[202]=77;
cos[203]=77;
cos[204]=77;
cos[205]=77;
cos[206]=77;
cos[207]=77;
cos[208]=77;
cos[209]=77;
cos[210]=77;
cos[211]=77;
cos[212]=77;
cos[213]=77;
cos[214]=77;
cos[215]=77;
cos[216]=77;
cos[217]=77;
cos[218]=77;
cos[219]=77;
cos[220]=77;
cos[221]=77;
cos[222]=77;
cos[223]=77;
cos[224]=77;
cos[225]=77;
cos[226]=77;
cos[227]=77;
cos[228]=77;
cos[229]=77;
cos[230]=77;
cos[231]=77;
cos[232]=77;
cos[233]=77;
cos[234]=77;
cos[235]=77;
cos[236]=77;
cos[237]=77;
cos[238]=77;
cos[239]=77;
cos[240]=77;
cos[241]=77;
cos[242]=77;
cos[243]=77;
cos[244]=77;
cos[245]=77;
cos[246]=77;
cos[247]=77;
cos[248]=77;
cos[249]=77;
cos[250]=77;
cos[251]=77;
cos[252]=77;
cos[253]=77;
cos[254]=77;
cos[255]=77;
cos[256]=77;
cos[257]=77;
cos[258]=77;
cos[259]=77;
cos[260]=77;
cos[261]=77;
cos[262]=77;
cos[263]=77;
cos[264]=77;
cos[265]=77;
cos[266]=77;
cos[267]=77;
cos[268]=77;
cos[269]=77;
cos[270]=77;
cos[271]=77;
cos[272]=77;
cos[273]=77;
cos[274]=77;
cos[275]=77;
cos[276]=77;
cos[277]=77;
cos[278]=77;
cos[279]=77;
cos[280]=77;
cos[281]=77;
cos[282]=77;
cos[283]=77;
cos[284]=77;
cos[285]=77;
cos[286]=77;
cos[287]=77;
cos[288]=77;
cos[289]=77;
cos[290]=77;
cos[291]=77;
cos[292]=77;
cos[293]=77;
cos[294]=77;
cos[295]=77;
cos[296]=77;
cos[297]=77;
cos[298]=77;
cos[299]=77;
cos[300]=77;
cos[301]=77;
cos[302]=77;
cos[303]=77;
cos[304]=77;
cos[305]=77;
cos[306]=77;
cos[307]=77;
cos[308]=77;
cos[309]=77;
cos[310]=77;
cos[311]=77;
cos[312]=77;
cos[313]=77;
cos[314]=77;
cos[315]=77;
cos[316]=77;
cos[317]=77;
cos[318]=77;
cos[319]=77;
cos[320]=77;
cos[321]=77;
cos[322]=77;
cos[323]=77;
cos[324]=77;
cos[325]=77;
cos[326]=76;
cos[327]=76;
cos[328]=76;
cos[329]=76;
cos[330]=76;
cos[331]=76;
cos[332]=76;
cos[333]=76;
cos[334]=76;
cos[335]=76;
cos[336]=76;
cos[337]=76;
cos[338]=76;
cos[339]=76;
cos[340]=76;
cos[341]=76;
cos[342]=76;
cos[343]=76;
cos[344]=76;
cos[345]=76;
cos[346]=76;
cos[347]=76;
cos[348]=76;
cos[349]=76;
cos[350]=76;
cos[351]=76;
cos[352]=76;
cos[353]=76;
cos[354]=76;
cos[355]=76;
cos[356]=76;
cos[357]=76;
cos[358]=76;
cos[359]=76;
cos[360]=76;
cos[361]=76;
cos[362]=76;
cos[363]=76;
cos[364]=76;
cos[365]=76;
cos[366]=76;
cos[367]=76;
cos[368]=76;
cos[369]=76;
cos[370]=76;
cos[371]=76;
cos[372]=76;
cos[373]=76;
cos[374]=76;
cos[375]=76;
cos[376]=76;
cos[377]=76;
cos[378]=76;
cos[379]=76;
cos[380]=76;
cos[381]=76;
cos[382]=76;
cos[383]=76;
cos[384]=76;
cos[385]=76;
cos[386]=76;
cos[387]=76;
cos[388]=76;
cos[389]=76;
cos[390]=76;
cos[391]=76;
cos[392]=76;
cos[393]=76;
cos[394]=76;
cos[395]=76;
cos[396]=76;
cos[397]=76;
cos[398]=76;
cos[399]=76;
cos[400]=76;
cos[401]=76;
cos[402]=76;
cos[403]=76;
cos[404]=76;
cos[405]=76;
cos[406]=76;
cos[407]=76;
cos[408]=76;
cos[409]=76;
cos[410]=76;
cos[411]=76;
cos[412]=76;
cos[413]=76;
cos[414]=75;
cos[415]=75;
cos[416]=75;
cos[417]=75;
cos[418]=75;
cos[419]=75;
cos[420]=75;
cos[421]=75;
cos[422]=75;
cos[423]=75;
cos[424]=75;
cos[425]=75;
cos[426]=75;
cos[427]=75;
cos[428]=75;
cos[429]=75;
cos[430]=75;
cos[431]=75;
cos[432]=75;
cos[433]=75;
cos[434]=75;
cos[435]=75;
cos[436]=75;
cos[437]=75;
cos[438]=75;
cos[439]=75;
cos[440]=75;
cos[441]=75;
cos[442]=75;
cos[443]=75;
cos[444]=75;
cos[445]=75;
cos[446]=75;
cos[447]=75;
cos[448]=75;
cos[449]=75;
cos[450]=75;
cos[451]=75;
cos[452]=75;
cos[453]=75;
cos[454]=75;
cos[455]=75;
cos[456]=75;
cos[457]=75;
cos[458]=75;
cos[459]=75;
cos[460]=75;
cos[461]=75;
cos[462]=75;
cos[463]=75;
cos[464]=75;
cos[465]=75;
cos[466]=75;
cos[467]=75;
cos[468]=75;
cos[469]=75;
cos[470]=75;
cos[471]=75;
cos[472]=75;
cos[473]=75;
cos[474]=75;
cos[475]=75;
cos[476]=75;
cos[477]=75;
cos[478]=75;
cos[479]=75;
cos[480]=75;
cos[481]=75;
cos[482]=75;
cos[483]=75;
cos[484]=75;
cos[485]=75;
cos[486]=75;
cos[487]=74;
cos[488]=74;
cos[489]=74;
cos[490]=74;
cos[491]=74;
cos[492]=74;
cos[493]=74;
cos[494]=74;
cos[495]=74;
cos[496]=74;
cos[497]=74;
cos[498]=74;
cos[499]=74;
cos[500]=74;
cos[501]=74;
cos[502]=74;
cos[503]=74;
cos[504]=74;
cos[505]=74;
cos[506]=74;
cos[507]=74;
cos[508]=74;
cos[509]=74;
cos[510]=74;
cos[511]=74;
cos[512]=74;
cos[513]=74;
cos[514]=74;
cos[515]=74;
cos[516]=74;
cos[517]=74;
cos[518]=74;
cos[519]=74;
cos[520]=74;
cos[521]=74;
cos[522]=74;
cos[523]=74;
cos[524]=74;
cos[525]=74;
cos[526]=74;
cos[527]=74;
cos[528]=74;
cos[529]=74;
cos[530]=74;
cos[531]=74;
cos[532]=74;
cos[533]=74;
cos[534]=74;
cos[535]=74;
cos[536]=74;
cos[537]=74;
cos[538]=74;
cos[539]=74;
cos[540]=74;
cos[541]=74;
cos[542]=74;
cos[543]=74;
cos[544]=74;
cos[545]=74;
cos[546]=74;
cos[547]=74;
cos[548]=74;
cos[549]=74;
cos[550]=74;
cos[551]=73;
cos[552]=73;
cos[553]=73;
cos[554]=73;
cos[555]=73;
cos[556]=73;
cos[557]=73;
cos[558]=73;
cos[559]=73;
cos[560]=73;
cos[561]=73;
cos[562]=73;
cos[563]=73;
cos[564]=73;
cos[565]=73;
cos[566]=73;
cos[567]=73;
cos[568]=73;
cos[569]=73;
cos[570]=73;
cos[571]=73;
cos[572]=73;
cos[573]=73;
cos[574]=73;
cos[575]=73;
cos[576]=73;
cos[577]=73;
cos[578]=73;
cos[579]=73;
cos[580]=73;
cos[581]=73;
cos[582]=73;
cos[583]=73;
cos[584]=73;
cos[585]=73;
cos[586]=73;
cos[587]=73;
cos[588]=73;
cos[589]=73;
cos[590]=73;
cos[591]=73;
cos[592]=73;
cos[593]=73;
cos[594]=73;
cos[595]=73;
cos[596]=73;
cos[597]=73;
cos[598]=73;
cos[599]=73;
cos[600]=73;
cos[601]=73;
cos[602]=73;
cos[603]=73;
cos[604]=73;
cos[605]=73;
cos[606]=73;
cos[607]=73;
cos[608]=72;
cos[609]=72;
cos[610]=72;
cos[611]=72;
cos[612]=72;
cos[613]=72;
cos[614]=72;
cos[615]=72;
cos[616]=72;
cos[617]=72;
cos[618]=72;
cos[619]=72;
cos[620]=72;
cos[621]=72;
cos[622]=72;
cos[623]=72;
cos[624]=72;
cos[625]=72;
cos[626]=72;
cos[627]=72;
cos[628]=72;
cos[629]=72;
cos[630]=72;
cos[631]=72;
cos[632]=72;
cos[633]=72;
cos[634]=72;
cos[635]=72;
cos[636]=72;
cos[637]=72;
cos[638]=72;
cos[639]=72;
cos[640]=72;
cos[641]=72;
cos[642]=72;
cos[643]=72;
cos[644]=72;
cos[645]=72;
cos[646]=72;
cos[647]=72;
cos[648]=72;
cos[649]=72;
cos[650]=72;
cos[651]=72;
cos[652]=72;
cos[653]=72;
cos[654]=72;
cos[655]=72;
cos[656]=72;
cos[657]=72;
cos[658]=72;
cos[659]=72;
cos[660]=72;
cos[661]=71;
cos[662]=71;
cos[663]=71;
cos[664]=71;
cos[665]=71;
cos[666]=71;
cos[667]=71;
cos[668]=71;
cos[669]=71;
cos[670]=71;
cos[671]=71;
cos[672]=71;
cos[673]=71;
cos[674]=71;
cos[675]=71;
cos[676]=71;
cos[677]=71;
cos[678]=71;
cos[679]=71;
cos[680]=71;
cos[681]=71;
cos[682]=71;
cos[683]=71;
cos[684]=71;
cos[685]=71;
cos[686]=71;
cos[687]=71;
cos[688]=71;
cos[689]=71;
cos[690]=71;
cos[691]=71;
cos[692]=71;
cos[693]=71;
cos[694]=71;
cos[695]=71;
cos[696]=71;
cos[697]=71;
cos[698]=71;
cos[699]=71;
cos[700]=71;
cos[701]=71;
cos[702]=71;
cos[703]=71;
cos[704]=71;
cos[705]=71;
cos[706]=71;
cos[707]=71;
cos[708]=71;
cos[709]=71;
cos[710]=70;
cos[711]=70;
cos[712]=70;
cos[713]=70;
cos[714]=70;
cos[715]=70;
cos[716]=70;
cos[717]=70;
cos[718]=70;
cos[719]=70;
cos[720]=70;
cos[721]=70;
cos[722]=70;
cos[723]=70;
cos[724]=70;
cos[725]=70;
cos[726]=70;
cos[727]=70;
cos[728]=70;
cos[729]=70;
cos[730]=70;
cos[731]=70;
cos[732]=70;
cos[733]=70;
cos[734]=70;
cos[735]=70;
cos[736]=70;
cos[737]=70;
cos[738]=70;
cos[739]=70;
cos[740]=70;
cos[741]=70;
cos[742]=70;
cos[743]=70;
cos[744]=70;
cos[745]=70;
cos[746]=70;
cos[747]=70;
cos[748]=70;
cos[749]=70;
cos[750]=70;
cos[751]=70;
cos[752]=70;
cos[753]=70;
cos[754]=70;
cos[755]=69;
cos[756]=69;
cos[757]=69;
cos[758]=69;
cos[759]=69;
cos[760]=69;
cos[761]=69;
cos[762]=69;
cos[763]=69;
cos[764]=69;
cos[765]=69;
cos[766]=69;
cos[767]=69;
cos[768]=69;
cos[769]=69;
cos[770]=69;
cos[771]=69;
cos[772]=69;
cos[773]=69;
cos[774]=69;
cos[775]=69;
cos[776]=69;
cos[777]=69;
cos[778]=69;
cos[779]=69;
cos[780]=69;
cos[781]=69;
cos[782]=69;
cos[783]=69;
cos[784]=69;
cos[785]=69;
cos[786]=69;
cos[787]=69;
cos[788]=69;
cos[789]=69;
cos[790]=69;
cos[791]=69;
cos[792]=69;
cos[793]=69;
cos[794]=69;
cos[795]=69;
cos[796]=69;
cos[797]=69;
cos[798]=69;
cos[799]=68;
cos[800]=68;
cos[801]=68;
cos[802]=68;
cos[803]=68;
cos[804]=68;
cos[805]=68;
cos[806]=68;
cos[807]=68;
cos[808]=68;
cos[809]=68;
cos[810]=68;
cos[811]=68;
cos[812]=68;
cos[813]=68;
cos[814]=68;
cos[815]=68;
cos[816]=68;
cos[817]=68;
cos[818]=68;
cos[819]=68;
cos[820]=68;
cos[821]=68;
cos[822]=68;
cos[823]=68;
cos[824]=68;
cos[825]=68;
cos[826]=68;
cos[827]=68;
cos[828]=68;
cos[829]=68;
cos[830]=68;
cos[831]=68;
cos[832]=68;
cos[833]=68;
cos[834]=68;
cos[835]=68;
cos[836]=68;
cos[837]=68;
cos[838]=68;
cos[839]=68;
cos[840]=67;
cos[841]=67;
cos[842]=67;
cos[843]=67;
cos[844]=67;
cos[845]=67;
cos[846]=67;
cos[847]=67;
cos[848]=67;
cos[849]=67;
cos[850]=67;
cos[851]=67;
cos[852]=67;
cos[853]=67;
cos[854]=67;
cos[855]=67;
cos[856]=67;
cos[857]=67;
cos[858]=67;
cos[859]=67;
cos[860]=67;
cos[861]=67;
cos[862]=67;
cos[863]=67;
cos[864]=67;
cos[865]=67;
cos[866]=67;
cos[867]=67;
cos[868]=67;
cos[869]=67;
cos[870]=67;
cos[871]=67;
cos[872]=67;
cos[873]=67;
cos[874]=67;
cos[875]=67;
cos[876]=67;
cos[877]=67;
cos[878]=67;
cos[879]=67;
cos[880]=66;
cos[881]=66;
cos[882]=66;
cos[883]=66;
cos[884]=66;
cos[885]=66;
cos[886]=66;
cos[887]=66;
cos[888]=66;
cos[889]=66;
cos[890]=66;
cos[891]=66;
cos[892]=66;
cos[893]=66;
cos[894]=66;
cos[895]=66;
cos[896]=66;
cos[897]=66;
cos[898]=66;
cos[899]=66;
cos[900]=66;
cos[901]=66;
cos[902]=66;
cos[903]=66;
cos[904]=66;
cos[905]=66;
cos[906]=66;
cos[907]=66;
cos[908]=66;
cos[909]=66;
cos[910]=66;
cos[911]=66;
cos[912]=66;
cos[913]=66;
cos[914]=66;
cos[915]=66;
cos[916]=66;
cos[917]=66;
cos[918]=65;
cos[919]=65;
cos[920]=65;
cos[921]=65;
cos[922]=65;
cos[923]=65;
cos[924]=65;
cos[925]=65;
cos[926]=65;
cos[927]=65;
cos[928]=65;
cos[929]=65;
cos[930]=65;
cos[931]=65;
cos[932]=65;
cos[933]=65;
cos[934]=65;
cos[935]=65;
cos[936]=65;
cos[937]=65;
cos[938]=65;
cos[939]=65;
cos[940]=65;
cos[941]=65;
cos[942]=65;
cos[943]=65;
cos[944]=65;
cos[945]=65;
cos[946]=65;
cos[947]=65;
cos[948]=65;
cos[949]=65;
cos[950]=65;
cos[951]=65;
cos[952]=65;
cos[953]=65;
cos[954]=65;
cos[955]=64;
cos[956]=64;
cos[957]=64;
cos[958]=64;
cos[959]=64;
cos[960]=64;
cos[961]=64;
cos[962]=64;
cos[963]=64;
cos[964]=64;
cos[965]=64;
cos[966]=64;
cos[967]=64;
cos[968]=64;
cos[969]=64;
cos[970]=64;
cos[971]=64;
cos[972]=64;
cos[973]=64;
cos[974]=64;
cos[975]=64;
cos[976]=64;
cos[977]=64;
cos[978]=64;
cos[979]=64;
cos[980]=64;
cos[981]=64;
cos[982]=64;
cos[983]=64;
cos[984]=64;
cos[985]=64;
cos[986]=64;
cos[987]=64;
cos[988]=64;
cos[989]=64;
cos[990]=63;
cos[991]=63;
cos[992]=63;
cos[993]=63;
cos[994]=63;
cos[995]=63;
cos[996]=63;
cos[997]=63;
cos[998]=63;
cos[999]=63;
cos[1000]=63;
cos[1001]=63;
cos[1002]=63;
cos[1003]=63;
cos[1004]=63;
cos[1005]=63;
cos[1006]=63;
cos[1007]=63;
cos[1008]=63;
cos[1009]=63;
cos[1010]=63;
cos[1011]=63;
cos[1012]=63;
cos[1013]=63;
cos[1014]=63;
cos[1015]=63;
cos[1016]=63;
cos[1017]=63;
cos[1018]=63;
cos[1019]=63;
cos[1020]=63;
cos[1021]=63;
cos[1022]=63;
cos[1023]=63;
cos[1024]=63;
cos[1025]=62;
cos[1026]=62;
cos[1027]=62;
cos[1028]=62;
cos[1029]=62;
cos[1030]=62;
cos[1031]=62;
cos[1032]=62;
cos[1033]=62;
cos[1034]=62;
cos[1035]=62;
cos[1036]=62;
cos[1037]=62;
cos[1038]=62;
cos[1039]=62;
cos[1040]=62;
cos[1041]=62;
cos[1042]=62;
cos[1043]=62;
cos[1044]=62;
cos[1045]=62;
cos[1046]=62;
cos[1047]=62;
cos[1048]=62;
cos[1049]=62;
cos[1050]=62;
cos[1051]=62;
cos[1052]=62;
cos[1053]=62;
cos[1054]=62;
cos[1055]=62;
cos[1056]=62;
cos[1057]=62;
cos[1058]=61;
cos[1059]=61;
cos[1060]=61;
cos[1061]=61;
cos[1062]=61;
cos[1063]=61;
cos[1064]=61;
cos[1065]=61;
cos[1066]=61;
cos[1067]=61;
cos[1068]=61;
cos[1069]=61;
cos[1070]=61;
cos[1071]=61;
cos[1072]=61;
cos[1073]=61;
cos[1074]=61;
cos[1075]=61;
cos[1076]=61;
cos[1077]=61;
cos[1078]=61;
cos[1079]=61;
cos[1080]=61;
cos[1081]=61;
cos[1082]=61;
cos[1083]=61;
cos[1084]=61;
cos[1085]=61;
cos[1086]=61;
cos[1087]=61;
cos[1088]=61;
cos[1089]=61;
cos[1090]=61;
cos[1091]=60;
cos[1092]=60;
cos[1093]=60;
cos[1094]=60;
cos[1095]=60;
cos[1096]=60;
cos[1097]=60;
cos[1098]=60;
cos[1099]=60;
cos[1100]=60;
cos[1101]=60;
cos[1102]=60;
cos[1103]=60;
cos[1104]=60;
cos[1105]=60;
cos[1106]=60;
cos[1107]=60;
cos[1108]=60;
cos[1109]=60;
cos[1110]=60;
cos[1111]=60;
cos[1112]=60;
cos[1113]=60;
cos[1114]=60;
cos[1115]=60;
cos[1116]=60;
cos[1117]=60;
cos[1118]=60;
cos[1119]=60;
cos[1120]=60;
cos[1121]=60;
cos[1122]=60;
cos[1123]=59;
cos[1124]=59;
cos[1125]=59;
cos[1126]=59;
cos[1127]=59;
cos[1128]=59;
cos[1129]=59;
cos[1130]=59;
cos[1131]=59;
cos[1132]=59;
cos[1133]=59;
cos[1134]=59;
cos[1135]=59;
cos[1136]=59;
cos[1137]=59;
cos[1138]=59;
cos[1139]=59;
cos[1140]=59;
cos[1141]=59;
cos[1142]=59;
cos[1143]=59;
cos[1144]=59;
cos[1145]=59;
cos[1146]=59;
cos[1147]=59;
cos[1148]=59;
cos[1149]=59;
cos[1150]=59;
cos[1151]=59;
cos[1152]=59;
cos[1153]=59;
cos[1154]=58;
cos[1155]=58;
cos[1156]=58;
cos[1157]=58;
cos[1158]=58;
cos[1159]=58;
cos[1160]=58;
cos[1161]=58;
cos[1162]=58;
cos[1163]=58;
cos[1164]=58;
cos[1165]=58;
cos[1166]=58;
cos[1167]=58;
cos[1168]=58;
cos[1169]=58;
cos[1170]=58;
cos[1171]=58;
cos[1172]=58;
cos[1173]=58;
cos[1174]=58;
cos[1175]=58;
cos[1176]=58;
cos[1177]=58;
cos[1178]=58;
cos[1179]=58;
cos[1180]=58;
cos[1181]=58;
cos[1182]=58;
cos[1183]=58;
cos[1184]=57;
cos[1185]=57;
cos[1186]=57;
cos[1187]=57;
cos[1188]=57;
cos[1189]=57;
cos[1190]=57;
cos[1191]=57;
cos[1192]=57;
cos[1193]=57;
cos[1194]=57;
cos[1195]=57;
cos[1196]=57;
cos[1197]=57;
cos[1198]=57;
cos[1199]=57;
cos[1200]=57;
cos[1201]=57;
cos[1202]=57;
cos[1203]=57;
cos[1204]=57;
cos[1205]=57;
cos[1206]=57;
cos[1207]=57;
cos[1208]=57;
cos[1209]=57;
cos[1210]=57;
cos[1211]=57;
cos[1212]=57;
cos[1213]=57;
cos[1214]=56;
cos[1215]=56;
cos[1216]=56;
cos[1217]=56;
cos[1218]=56;
cos[1219]=56;
cos[1220]=56;
cos[1221]=56;
cos[1222]=56;
cos[1223]=56;
cos[1224]=56;
cos[1225]=56;
cos[1226]=56;
cos[1227]=56;
cos[1228]=56;
cos[1229]=56;
cos[1230]=56;
cos[1231]=56;
cos[1232]=56;
cos[1233]=56;
cos[1234]=56;
cos[1235]=56;
cos[1236]=56;
cos[1237]=56;
cos[1238]=56;
cos[1239]=56;
cos[1240]=56;
cos[1241]=56;
cos[1242]=56;
cos[1243]=55;
cos[1244]=55;
cos[1245]=55;
cos[1246]=55;
cos[1247]=55;
cos[1248]=55;
cos[1249]=55;
cos[1250]=55;
cos[1251]=55;
cos[1252]=55;
cos[1253]=55;
cos[1254]=55;
cos[1255]=55;
cos[1256]=55;
cos[1257]=55;
cos[1258]=55;
cos[1259]=55;
cos[1260]=55;
cos[1261]=55;
cos[1262]=55;
cos[1263]=55;
cos[1264]=55;
cos[1265]=55;
cos[1266]=55;
cos[1267]=55;
cos[1268]=55;
cos[1269]=55;
cos[1270]=55;
cos[1271]=55;
cos[1272]=54;
cos[1273]=54;
cos[1274]=54;
cos[1275]=54;
cos[1276]=54;
cos[1277]=54;
cos[1278]=54;
cos[1279]=54;
cos[1280]=54;
cos[1281]=54;
cos[1282]=54;
cos[1283]=54;
cos[1284]=54;
cos[1285]=54;
cos[1286]=54;
cos[1287]=54;
cos[1288]=54;
cos[1289]=54;
cos[1290]=54;
cos[1291]=54;
cos[1292]=54;
cos[1293]=54;
cos[1294]=54;
cos[1295]=54;
cos[1296]=54;
cos[1297]=54;
cos[1298]=54;
cos[1299]=54;
cos[1300]=53;
cos[1301]=53;
cos[1302]=53;
cos[1303]=53;
cos[1304]=53;
cos[1305]=53;
cos[1306]=53;
cos[1307]=53;
cos[1308]=53;
cos[1309]=53;
cos[1310]=53;
cos[1311]=53;
cos[1312]=53;
cos[1313]=53;
cos[1314]=53;
cos[1315]=53;
cos[1316]=53;
cos[1317]=53;
cos[1318]=53;
cos[1319]=53;
cos[1320]=53;
cos[1321]=53;
cos[1322]=53;
cos[1323]=53;
cos[1324]=53;
cos[1325]=53;
cos[1326]=53;
cos[1327]=53;
cos[1328]=52;
cos[1329]=52;
cos[1330]=52;
cos[1331]=52;
cos[1332]=52;
cos[1333]=52;
cos[1334]=52;
cos[1335]=52;
cos[1336]=52;
cos[1337]=52;
cos[1338]=52;
cos[1339]=52;
cos[1340]=52;
cos[1341]=52;
cos[1342]=52;
cos[1343]=52;
cos[1344]=52;
cos[1345]=52;
cos[1346]=52;
cos[1347]=52;
cos[1348]=52;
cos[1349]=52;
cos[1350]=52;
cos[1351]=52;
cos[1352]=52;
cos[1353]=52;
cos[1354]=52;
cos[1355]=51;
cos[1356]=51;
cos[1357]=51;
cos[1358]=51;
cos[1359]=51;
cos[1360]=51;
cos[1361]=51;
cos[1362]=51;
cos[1363]=51;
cos[1364]=51;
cos[1365]=51;
cos[1366]=51;
cos[1367]=51;
cos[1368]=51;
cos[1369]=51;
cos[1370]=51;
cos[1371]=51;
cos[1372]=51;
cos[1373]=51;
cos[1374]=51;
cos[1375]=51;
cos[1376]=51;
cos[1377]=51;
cos[1378]=51;
cos[1379]=51;
cos[1380]=51;
cos[1381]=51;
cos[1382]=50;
cos[1383]=50;
cos[1384]=50;
cos[1385]=50;
cos[1386]=50;
cos[1387]=50;
cos[1388]=50;
cos[1389]=50;
cos[1390]=50;
cos[1391]=50;
cos[1392]=50;
cos[1393]=50;
cos[1394]=50;
cos[1395]=50;
cos[1396]=50;
cos[1397]=50;
cos[1398]=50;
cos[1399]=50;
cos[1400]=50;
cos[1401]=50;
cos[1402]=50;
cos[1403]=50;
cos[1404]=50;
cos[1405]=50;
cos[1406]=50;
cos[1407]=50;
cos[1408]=49;
cos[1409]=49;
cos[1410]=49;
cos[1411]=49;
cos[1412]=49;
cos[1413]=49;
cos[1414]=49;
cos[1415]=49;
cos[1416]=49;
cos[1417]=49;
cos[1418]=49;
cos[1419]=49;
cos[1420]=49;
cos[1421]=49;
cos[1422]=49;
cos[1423]=49;
cos[1424]=49;
cos[1425]=49;
cos[1426]=49;
cos[1427]=49;
cos[1428]=49;
cos[1429]=49;
cos[1430]=49;
cos[1431]=49;
cos[1432]=49;
cos[1433]=49;
cos[1434]=49;
cos[1435]=48;
cos[1436]=48;
cos[1437]=48;
cos[1438]=48;
cos[1439]=48;
cos[1440]=48;
cos[1441]=48;
cos[1442]=48;
cos[1443]=48;
cos[1444]=48;
cos[1445]=48;
cos[1446]=48;
cos[1447]=48;
cos[1448]=48;
cos[1449]=48;
cos[1450]=48;
cos[1451]=48;
cos[1452]=48;
cos[1453]=48;
cos[1454]=48;
cos[1455]=48;
cos[1456]=48;
cos[1457]=48;
cos[1458]=48;
cos[1459]=48;
cos[1460]=47;
cos[1461]=47;
cos[1462]=47;
cos[1463]=47;
cos[1464]=47;
cos[1465]=47;
cos[1466]=47;
cos[1467]=47;
cos[1468]=47;
cos[1469]=47;
cos[1470]=47;
cos[1471]=47;
cos[1472]=47;
cos[1473]=47;
cos[1474]=47;
cos[1475]=47;
cos[1476]=47;
cos[1477]=47;
cos[1478]=47;
cos[1479]=47;
cos[1480]=47;
cos[1481]=47;
cos[1482]=47;
cos[1483]=47;
cos[1484]=47;
cos[1485]=47;
cos[1486]=46;
cos[1487]=46;
cos[1488]=46;
cos[1489]=46;
cos[1490]=46;
cos[1491]=46;
cos[1492]=46;
cos[1493]=46;
cos[1494]=46;
cos[1495]=46;
cos[1496]=46;
cos[1497]=46;
cos[1498]=46;
cos[1499]=46;
cos[1500]=46;
cos[1501]=46;
cos[1502]=46;
cos[1503]=46;
cos[1504]=46;
cos[1505]=46;
cos[1506]=46;
cos[1507]=46;
cos[1508]=46;
cos[1509]=46;
cos[1510]=46;
cos[1511]=45;
cos[1512]=45;
cos[1513]=45;
cos[1514]=45;
cos[1515]=45;
cos[1516]=45;
cos[1517]=45;
cos[1518]=45;
cos[1519]=45;
cos[1520]=45;
cos[1521]=45;
cos[1522]=45;
cos[1523]=45;
cos[1524]=45;
cos[1525]=45;
cos[1526]=45;
cos[1527]=45;
cos[1528]=45;
cos[1529]=45;
cos[1530]=45;
cos[1531]=45;
cos[1532]=45;
cos[1533]=45;
cos[1534]=45;
cos[1535]=45;
cos[1536]=44;
cos[1537]=44;
cos[1538]=44;
cos[1539]=44;
cos[1540]=44;
cos[1541]=44;
cos[1542]=44;
cos[1543]=44;
cos[1544]=44;
cos[1545]=44;
cos[1546]=44;
cos[1547]=44;
cos[1548]=44;
cos[1549]=44;
cos[1550]=44;
cos[1551]=44;
cos[1552]=44;
cos[1553]=44;
cos[1554]=44;
cos[1555]=44;
cos[1556]=44;
cos[1557]=44;
cos[1558]=44;
cos[1559]=44;
cos[1560]=44;
cos[1561]=43;
cos[1562]=43;
cos[1563]=43;
cos[1564]=43;
cos[1565]=43;
cos[1566]=43;
cos[1567]=43;
cos[1568]=43;
cos[1569]=43;
cos[1570]=43;
cos[1571]=43;
cos[1572]=43;
cos[1573]=43;
cos[1574]=43;
cos[1575]=43;
cos[1576]=43;
cos[1577]=43;
cos[1578]=43;
cos[1579]=43;
cos[1580]=43;
cos[1581]=43;
cos[1582]=43;
cos[1583]=43;
cos[1584]=43;
cos[1585]=42;
cos[1586]=42;
cos[1587]=42;
cos[1588]=42;
cos[1589]=42;
cos[1590]=42;
cos[1591]=42;
cos[1592]=42;
cos[1593]=42;
cos[1594]=42;
cos[1595]=42;
cos[1596]=42;
cos[1597]=42;
cos[1598]=42;
cos[1599]=42;
cos[1600]=42;
cos[1601]=42;
cos[1602]=42;
cos[1603]=42;
cos[1604]=42;
cos[1605]=42;
cos[1606]=42;
cos[1607]=42;
cos[1608]=42;
cos[1609]=41;
cos[1610]=41;
cos[1611]=41;
cos[1612]=41;
cos[1613]=41;
cos[1614]=41;
cos[1615]=41;
cos[1616]=41;
cos[1617]=41;
cos[1618]=41;
cos[1619]=41;
cos[1620]=41;
cos[1621]=41;
cos[1622]=41;
cos[1623]=41;
cos[1624]=41;
cos[1625]=41;
cos[1626]=41;
cos[1627]=41;
cos[1628]=41;
cos[1629]=41;
cos[1630]=41;
cos[1631]=41;
cos[1632]=41;
cos[1633]=40;
cos[1634]=40;
cos[1635]=40;
cos[1636]=40;
cos[1637]=40;
cos[1638]=40;
cos[1639]=40;
cos[1640]=40;
cos[1641]=40;
cos[1642]=40;
cos[1643]=40;
cos[1644]=40;
cos[1645]=40;
cos[1646]=40;
cos[1647]=40;
cos[1648]=40;
cos[1649]=40;
cos[1650]=40;
cos[1651]=40;
cos[1652]=40;
cos[1653]=40;
cos[1654]=40;
cos[1655]=40;
cos[1656]=40;
cos[1657]=39;
cos[1658]=39;
cos[1659]=39;
cos[1660]=39;
cos[1661]=39;
cos[1662]=39;
cos[1663]=39;
cos[1664]=39;
cos[1665]=39;
cos[1666]=39;
cos[1667]=39;
cos[1668]=39;
cos[1669]=39;
cos[1670]=39;
cos[1671]=39;
cos[1672]=39;
cos[1673]=39;
cos[1674]=39;
cos[1675]=39;
cos[1676]=39;
cos[1677]=39;
cos[1678]=39;
cos[1679]=39;
cos[1680]=38;
cos[1681]=38;
cos[1682]=38;
cos[1683]=38;
cos[1684]=38;
cos[1685]=38;
cos[1686]=38;
cos[1687]=38;
cos[1688]=38;
cos[1689]=38;
cos[1690]=38;
cos[1691]=38;
cos[1692]=38;
cos[1693]=38;
cos[1694]=38;
cos[1695]=38;
cos[1696]=38;
cos[1697]=38;
cos[1698]=38;
cos[1699]=38;
cos[1700]=38;
cos[1701]=38;
cos[1702]=38;
cos[1703]=38;
cos[1704]=37;
cos[1705]=37;
cos[1706]=37;
cos[1707]=37;
cos[1708]=37;
cos[1709]=37;
cos[1710]=37;
cos[1711]=37;
cos[1712]=37;
cos[1713]=37;
cos[1714]=37;
cos[1715]=37;
cos[1716]=37;
cos[1717]=37;
cos[1718]=37;
cos[1719]=37;
cos[1720]=37;
cos[1721]=37;
cos[1722]=37;
cos[1723]=37;
cos[1724]=37;
cos[1725]=37;
cos[1726]=37;
cos[1727]=36;
cos[1728]=36;
cos[1729]=36;
cos[1730]=36;
cos[1731]=36;
cos[1732]=36;
cos[1733]=36;
cos[1734]=36;
cos[1735]=36;
cos[1736]=36;
cos[1737]=36;
cos[1738]=36;
cos[1739]=36;
cos[1740]=36;
cos[1741]=36;
cos[1742]=36;
cos[1743]=36;
cos[1744]=36;
cos[1745]=36;
cos[1746]=36;
cos[1747]=36;
cos[1748]=36;
cos[1749]=36;
cos[1750]=35;
cos[1751]=35;
cos[1752]=35;
cos[1753]=35;
cos[1754]=35;
cos[1755]=35;
cos[1756]=35;
cos[1757]=35;
cos[1758]=35;
cos[1759]=35;
cos[1760]=35;
cos[1761]=35;
cos[1762]=35;
cos[1763]=35;
cos[1764]=35;
cos[1765]=35;
cos[1766]=35;
cos[1767]=35;
cos[1768]=35;
cos[1769]=35;
cos[1770]=35;
cos[1771]=35;
cos[1772]=35;
cos[1773]=34;
cos[1774]=34;
cos[1775]=34;
cos[1776]=34;
cos[1777]=34;
cos[1778]=34;
cos[1779]=34;
cos[1780]=34;
cos[1781]=34;
cos[1782]=34;
cos[1783]=34;
cos[1784]=34;
cos[1785]=34;
cos[1786]=34;
cos[1787]=34;
cos[1788]=34;
cos[1789]=34;
cos[1790]=34;
cos[1791]=34;
cos[1792]=34;
cos[1793]=34;
cos[1794]=34;
cos[1795]=33;
cos[1796]=33;
cos[1797]=33;
cos[1798]=33;
cos[1799]=33;
cos[1800]=33;
cos[1801]=33;
cos[1802]=33;
cos[1803]=33;
cos[1804]=33;
cos[1805]=33;
cos[1806]=33;
cos[1807]=33;
cos[1808]=33;
cos[1809]=33;
cos[1810]=33;
cos[1811]=33;
cos[1812]=33;
cos[1813]=33;
cos[1814]=33;
cos[1815]=33;
cos[1816]=33;
cos[1817]=33;
cos[1818]=32;
cos[1819]=32;
cos[1820]=32;
cos[1821]=32;
cos[1822]=32;
cos[1823]=32;
cos[1824]=32;
cos[1825]=32;
cos[1826]=32;
cos[1827]=32;
cos[1828]=32;
cos[1829]=32;
cos[1830]=32;
cos[1831]=32;
cos[1832]=32;
cos[1833]=32;
cos[1834]=32;
cos[1835]=32;
cos[1836]=32;
cos[1837]=32;
cos[1838]=32;
cos[1839]=32;
cos[1840]=31;
cos[1841]=31;
cos[1842]=31;
cos[1843]=31;
cos[1844]=31;
cos[1845]=31;
cos[1846]=31;
cos[1847]=31;
cos[1848]=31;
cos[1849]=31;
cos[1850]=31;
cos[1851]=31;
cos[1852]=31;
cos[1853]=31;
cos[1854]=31;
cos[1855]=31;
cos[1856]=31;
cos[1857]=31;
cos[1858]=31;
cos[1859]=31;
cos[1860]=31;
cos[1861]=31;
cos[1862]=30;
cos[1863]=30;
cos[1864]=30;
cos[1865]=30;
cos[1866]=30;
cos[1867]=30;
cos[1868]=30;
cos[1869]=30;
cos[1870]=30;
cos[1871]=30;
cos[1872]=30;
cos[1873]=30;
cos[1874]=30;
cos[1875]=30;
cos[1876]=30;
cos[1877]=30;
cos[1878]=30;
cos[1879]=30;
cos[1880]=30;
cos[1881]=30;
cos[1882]=30;
cos[1883]=30;
cos[1884]=29;
cos[1885]=29;
cos[1886]=29;
cos[1887]=29;
cos[1888]=29;
cos[1889]=29;
cos[1890]=29;
cos[1891]=29;
cos[1892]=29;
cos[1893]=29;
cos[1894]=29;
cos[1895]=29;
cos[1896]=29;
cos[1897]=29;
cos[1898]=29;
cos[1899]=29;
cos[1900]=29;
cos[1901]=29;
cos[1902]=29;
cos[1903]=29;
cos[1904]=29;
cos[1905]=29;
cos[1906]=28;
cos[1907]=28;
cos[1908]=28;
cos[1909]=28;
cos[1910]=28;
cos[1911]=28;
cos[1912]=28;
cos[1913]=28;
cos[1914]=28;
cos[1915]=28;
cos[1916]=28;
cos[1917]=28;
cos[1918]=28;
cos[1919]=28;
cos[1920]=28;
cos[1921]=28;
cos[1922]=28;
cos[1923]=28;
cos[1924]=28;
cos[1925]=28;
cos[1926]=28;
cos[1927]=28;
cos[1928]=27;
cos[1929]=27;
cos[1930]=27;
cos[1931]=27;
cos[1932]=27;
cos[1933]=27;
cos[1934]=27;
cos[1935]=27;
cos[1936]=27;
cos[1937]=27;
cos[1938]=27;
cos[1939]=27;
cos[1940]=27;
cos[1941]=27;
cos[1942]=27;
cos[1943]=27;
cos[1944]=27;
cos[1945]=27;
cos[1946]=27;
cos[1947]=27;
cos[1948]=27;
cos[1949]=27;
cos[1950]=26;
cos[1951]=26;
cos[1952]=26;
cos[1953]=26;
cos[1954]=26;
cos[1955]=26;
cos[1956]=26;
cos[1957]=26;
cos[1958]=26;
cos[1959]=26;
cos[1960]=26;
cos[1961]=26;
cos[1962]=26;
cos[1963]=26;
cos[1964]=26;
cos[1965]=26;
cos[1966]=26;
cos[1967]=26;
cos[1968]=26;
cos[1969]=26;
cos[1970]=26;
cos[1971]=25;
cos[1972]=25;
cos[1973]=25;
cos[1974]=25;
cos[1975]=25;
cos[1976]=25;
cos[1977]=25;
cos[1978]=25;
cos[1979]=25;
cos[1980]=25;
cos[1981]=25;
cos[1982]=25;
cos[1983]=25;
cos[1984]=25;
cos[1985]=25;
cos[1986]=25;
cos[1987]=25;
cos[1988]=25;
cos[1989]=25;
cos[1990]=25;
cos[1991]=25;
cos[1992]=25;
cos[1993]=24;
cos[1994]=24;
cos[1995]=24;
cos[1996]=24;
cos[1997]=24;
cos[1998]=24;
cos[1999]=24;
cos[2000]=24;
cos[2001]=24;
cos[2002]=24;
cos[2003]=24;
cos[2004]=24;
cos[2005]=24;
cos[2006]=24;
cos[2007]=24;
cos[2008]=24;
cos[2009]=24;
cos[2010]=24;
cos[2011]=24;
cos[2012]=24;
cos[2013]=24;
cos[2014]=23;
cos[2015]=23;
cos[2016]=23;
cos[2017]=23;
cos[2018]=23;
cos[2019]=23;
cos[2020]=23;
cos[2021]=23;
cos[2022]=23;
cos[2023]=23;
cos[2024]=23;
cos[2025]=23;
cos[2026]=23;
cos[2027]=23;
cos[2028]=23;
cos[2029]=23;
cos[2030]=23;
cos[2031]=23;
cos[2032]=23;
cos[2033]=23;
cos[2034]=23;
cos[2035]=23;
cos[2036]=22;
cos[2037]=22;
cos[2038]=22;
cos[2039]=22;
cos[2040]=22;
cos[2041]=22;
cos[2042]=22;
cos[2043]=22;
cos[2044]=22;
cos[2045]=22;
cos[2046]=22;
cos[2047]=22;
cos[2048]=22;
cos[2049]=22;
cos[2050]=22;
cos[2051]=22;
cos[2052]=22;
cos[2053]=22;
cos[2054]=22;
cos[2055]=22;
cos[2056]=22;
cos[2057]=21;
cos[2058]=21;
cos[2059]=21;
cos[2060]=21;
cos[2061]=21;
cos[2062]=21;
cos[2063]=21;
cos[2064]=21;
cos[2065]=21;
cos[2066]=21;
cos[2067]=21;
cos[2068]=21;
cos[2069]=21;
cos[2070]=21;
cos[2071]=21;
cos[2072]=21;
cos[2073]=21;
cos[2074]=21;
cos[2075]=21;
cos[2076]=21;
cos[2077]=21;
cos[2078]=20;
cos[2079]=20;
cos[2080]=20;
cos[2081]=20;
cos[2082]=20;
cos[2083]=20;
cos[2084]=20;
cos[2085]=20;
cos[2086]=20;
cos[2087]=20;
cos[2088]=20;
cos[2089]=20;
cos[2090]=20;
cos[2091]=20;
cos[2092]=20;
cos[2093]=20;
cos[2094]=20;
cos[2095]=20;
cos[2096]=20;
cos[2097]=20;
cos[2098]=20;
cos[2099]=19;
cos[2100]=19;
cos[2101]=19;
cos[2102]=19;
cos[2103]=19;
cos[2104]=19;
cos[2105]=19;
cos[2106]=19;
cos[2107]=19;
cos[2108]=19;
cos[2109]=19;
cos[2110]=19;
cos[2111]=19;
cos[2112]=19;
cos[2113]=19;
cos[2114]=19;
cos[2115]=19;
cos[2116]=19;
cos[2117]=19;
cos[2118]=19;
cos[2119]=19;
cos[2120]=18;
cos[2121]=18;
cos[2122]=18;
cos[2123]=18;
cos[2124]=18;
cos[2125]=18;
cos[2126]=18;
cos[2127]=18;
cos[2128]=18;
cos[2129]=18;
cos[2130]=18;
cos[2131]=18;
cos[2132]=18;
cos[2133]=18;
cos[2134]=18;
cos[2135]=18;
cos[2136]=18;
cos[2137]=18;
cos[2138]=18;
cos[2139]=18;
cos[2140]=18;
cos[2141]=17;
cos[2142]=17;
cos[2143]=17;
cos[2144]=17;
cos[2145]=17;
cos[2146]=17;
cos[2147]=17;
cos[2148]=17;
cos[2149]=17;
cos[2150]=17;
cos[2151]=17;
cos[2152]=17;
cos[2153]=17;
cos[2154]=17;
cos[2155]=17;
cos[2156]=17;
cos[2157]=17;
cos[2158]=17;
cos[2159]=17;
cos[2160]=17;
cos[2161]=17;
cos[2162]=16;
cos[2163]=16;
cos[2164]=16;
cos[2165]=16;
cos[2166]=16;
cos[2167]=16;
cos[2168]=16;
cos[2169]=16;
cos[2170]=16;
cos[2171]=16;
cos[2172]=16;
cos[2173]=16;
cos[2174]=16;
cos[2175]=16;
cos[2176]=16;
cos[2177]=16;
cos[2178]=16;
cos[2179]=16;
cos[2180]=16;
cos[2181]=16;
cos[2182]=16;
cos[2183]=15;
cos[2184]=15;
cos[2185]=15;
cos[2186]=15;
cos[2187]=15;
cos[2188]=15;
cos[2189]=15;
cos[2190]=15;
cos[2191]=15;
cos[2192]=15;
cos[2193]=15;
cos[2194]=15;
cos[2195]=15;
cos[2196]=15;
cos[2197]=15;
cos[2198]=15;
cos[2199]=15;
cos[2200]=15;
cos[2201]=15;
cos[2202]=15;
cos[2203]=14;
cos[2204]=14;
cos[2205]=14;
cos[2206]=14;
cos[2207]=14;
cos[2208]=14;
cos[2209]=14;
cos[2210]=14;
cos[2211]=14;
cos[2212]=14;
cos[2213]=14;
cos[2214]=14;
cos[2215]=14;
cos[2216]=14;
cos[2217]=14;
cos[2218]=14;
cos[2219]=14;
cos[2220]=14;
cos[2221]=14;
cos[2222]=14;
cos[2223]=14;
cos[2224]=13;
cos[2225]=13;
cos[2226]=13;
cos[2227]=13;
cos[2228]=13;
cos[2229]=13;
cos[2230]=13;
cos[2231]=13;
cos[2232]=13;
cos[2233]=13;
cos[2234]=13;
cos[2235]=13;
cos[2236]=13;
cos[2237]=13;
cos[2238]=13;
cos[2239]=13;
cos[2240]=13;
cos[2241]=13;
cos[2242]=13;
cos[2243]=13;
cos[2244]=13;
cos[2245]=12;
cos[2246]=12;
cos[2247]=12;
cos[2248]=12;
cos[2249]=12;
cos[2250]=12;
cos[2251]=12;
cos[2252]=12;
cos[2253]=12;
cos[2254]=12;
cos[2255]=12;
cos[2256]=12;
cos[2257]=12;
cos[2258]=12;
cos[2259]=12;
cos[2260]=12;
cos[2261]=12;
cos[2262]=12;
cos[2263]=12;
cos[2264]=12;
cos[2265]=11;
cos[2266]=11;
cos[2267]=11;
cos[2268]=11;
cos[2269]=11;
cos[2270]=11;
cos[2271]=11;
cos[2272]=11;
cos[2273]=11;
cos[2274]=11;
cos[2275]=11;
cos[2276]=11;
cos[2277]=11;
cos[2278]=11;
cos[2279]=11;
cos[2280]=11;
cos[2281]=11;
cos[2282]=11;
cos[2283]=11;
cos[2284]=11;
cos[2285]=11;
cos[2286]=10;
cos[2287]=10;
cos[2288]=10;
cos[2289]=10;
cos[2290]=10;
cos[2291]=10;
cos[2292]=10;
cos[2293]=10;
cos[2294]=10;
cos[2295]=10;
cos[2296]=10;
cos[2297]=10;
cos[2298]=10;
cos[2299]=10;
cos[2300]=10;
cos[2301]=10;
cos[2302]=10;
cos[2303]=10;
cos[2304]=10;
cos[2305]=10;
cos[2306]=9;
cos[2307]=9;
cos[2308]=9;
cos[2309]=9;
cos[2310]=9;
cos[2311]=9;
cos[2312]=9;
cos[2313]=9;
cos[2314]=9;
cos[2315]=9;
cos[2316]=9;
cos[2317]=9;
cos[2318]=9;
cos[2319]=9;
cos[2320]=9;
cos[2321]=9;
cos[2322]=9;
cos[2323]=9;
cos[2324]=9;
cos[2325]=9;
cos[2326]=9;
cos[2327]=8;
cos[2328]=8;
cos[2329]=8;
cos[2330]=8;
cos[2331]=8;
cos[2332]=8;
cos[2333]=8;
cos[2334]=8;
cos[2335]=8;
cos[2336]=8;
cos[2337]=8;
cos[2338]=8;
cos[2339]=8;
cos[2340]=8;
cos[2341]=8;
cos[2342]=8;
cos[2343]=8;
cos[2344]=8;
cos[2345]=8;
cos[2346]=8;
cos[2347]=7;
cos[2348]=7;
cos[2349]=7;
cos[2350]=7;
cos[2351]=7;
cos[2352]=7;
cos[2353]=7;
cos[2354]=7;
cos[2355]=7;
cos[2356]=7;
cos[2357]=7;
cos[2358]=7;
cos[2359]=7;
cos[2360]=7;
cos[2361]=7;
cos[2362]=7;
cos[2363]=7;
cos[2364]=7;
cos[2365]=7;
cos[2366]=7;
cos[2367]=7;
cos[2368]=6;
cos[2369]=6;
cos[2370]=6;
cos[2371]=6;
cos[2372]=6;
cos[2373]=6;
cos[2374]=6;
cos[2375]=6;
cos[2376]=6;
cos[2377]=6;
cos[2378]=6;
cos[2379]=6;
cos[2380]=6;
cos[2381]=6;
cos[2382]=6;
cos[2383]=6;
cos[2384]=6;
cos[2385]=6;
cos[2386]=6;
cos[2387]=6;
cos[2388]=5;
cos[2389]=5;
cos[2390]=5;
cos[2391]=5;
cos[2392]=5;
cos[2393]=5;
cos[2394]=5;
cos[2395]=5;
cos[2396]=5;
cos[2397]=5;
cos[2398]=5;
cos[2399]=5;
cos[2400]=5;
cos[2401]=5;
cos[2402]=5;
cos[2403]=5;
cos[2404]=5;
cos[2405]=5;
cos[2406]=5;
cos[2407]=5;
cos[2408]=5;
cos[2409]=4;
cos[2410]=4;
cos[2411]=4;
cos[2412]=4;
cos[2413]=4;
cos[2414]=4;
cos[2415]=4;
cos[2416]=4;
cos[2417]=4;
cos[2418]=4;
cos[2419]=4;
cos[2420]=4;
cos[2421]=4;
cos[2422]=4;
cos[2423]=4;
cos[2424]=4;
cos[2425]=4;
cos[2426]=4;
cos[2427]=4;
cos[2428]=4;
cos[2429]=3;
cos[2430]=3;
cos[2431]=3;
cos[2432]=3;
cos[2433]=3;
cos[2434]=3;
cos[2435]=3;
cos[2436]=3;
cos[2437]=3;
cos[2438]=3;
cos[2439]=3;
cos[2440]=3;
cos[2441]=3;
cos[2442]=3;
cos[2443]=3;
cos[2444]=3;
cos[2445]=3;
cos[2446]=3;
cos[2447]=3;
cos[2448]=3;
cos[2449]=3;
cos[2450]=2;
cos[2451]=2;
cos[2452]=2;
cos[2453]=2;
cos[2454]=2;
cos[2455]=2;
cos[2456]=2;
cos[2457]=2;
cos[2458]=2;
cos[2459]=2;
cos[2460]=2;
cos[2461]=2;
cos[2462]=2;
cos[2463]=2;
cos[2464]=2;
cos[2465]=2;
cos[2466]=2;
cos[2467]=2;
cos[2468]=2;
cos[2469]=2;
cos[2470]=1;
cos[2471]=1;
cos[2472]=1;
cos[2473]=1;
cos[2474]=1;
cos[2475]=1;
cos[2476]=1;
cos[2477]=1;
cos[2478]=1;
cos[2479]=1;
cos[2480]=1;
cos[2481]=1;
cos[2482]=1;
cos[2483]=1;
cos[2484]=1;
cos[2485]=1;
cos[2486]=1;
cos[2487]=1;
cos[2488]=1;
cos[2489]=1;
cos[2490]=0;
cos[2491]=0;
cos[2492]=0;
cos[2493]=0;
cos[2494]=0;
cos[2495]=0;
cos[2496]=0;
cos[2497]=0;
cos[2498]=0;
cos[2499]=0;
cos[2500]=0;
cos[2501]=0;
cos[2502]=0;
cos[2503]=0;
cos[2504]=0;
cos[2505]=0;
cos[2506]=0;
cos[2507]=0;
cos[2508]=0;
cos[2509]=0;
cos[2510]=0;
cos[2511]=-1;
cos[2512]=-1;
cos[2513]=-1;
cos[2514]=-1;
cos[2515]=-1;
cos[2516]=-1;
cos[2517]=-1;
cos[2518]=-1;
cos[2519]=-1;
cos[2520]=-1;
cos[2521]=-1;
cos[2522]=-1;
cos[2523]=-1;
cos[2524]=-1;
cos[2525]=-1;
cos[2526]=-1;
cos[2527]=-1;
cos[2528]=-1;
cos[2529]=-1;
cos[2530]=-1;
cos[2531]=-2;
cos[2532]=-2;
cos[2533]=-2;
cos[2534]=-2;
cos[2535]=-2;
cos[2536]=-2;
cos[2537]=-2;
cos[2538]=-2;
cos[2539]=-2;
cos[2540]=-2;
cos[2541]=-2;
cos[2542]=-2;
cos[2543]=-2;
cos[2544]=-2;
cos[2545]=-2;
cos[2546]=-2;
cos[2547]=-2;
cos[2548]=-2;
cos[2549]=-2;
cos[2550]=-2;
cos[2551]=-3;
cos[2552]=-3;
cos[2553]=-3;
cos[2554]=-3;
cos[2555]=-3;
cos[2556]=-3;
cos[2557]=-3;
cos[2558]=-3;
cos[2559]=-3;
cos[2560]=-3;
cos[2561]=-3;
cos[2562]=-3;
cos[2563]=-3;
cos[2564]=-3;
cos[2565]=-3;
cos[2566]=-3;
cos[2567]=-3;
cos[2568]=-3;
cos[2569]=-3;
cos[2570]=-3;
cos[2571]=-3;
cos[2572]=-4;
cos[2573]=-4;
cos[2574]=-4;
cos[2575]=-4;
cos[2576]=-4;
cos[2577]=-4;
cos[2578]=-4;
cos[2579]=-4;
cos[2580]=-4;
cos[2581]=-4;
cos[2582]=-4;
cos[2583]=-4;
cos[2584]=-4;
cos[2585]=-4;
cos[2586]=-4;
cos[2587]=-4;
cos[2588]=-4;
cos[2589]=-4;
cos[2590]=-4;
cos[2591]=-4;
cos[2592]=-5;
cos[2593]=-5;
cos[2594]=-5;
cos[2595]=-5;
cos[2596]=-5;
cos[2597]=-5;
cos[2598]=-5;
cos[2599]=-5;
cos[2600]=-5;
cos[2601]=-5;
cos[2602]=-5;
cos[2603]=-5;
cos[2604]=-5;
cos[2605]=-5;
cos[2606]=-5;
cos[2607]=-5;
cos[2608]=-5;
cos[2609]=-5;
cos[2610]=-5;
cos[2611]=-5;
cos[2612]=-5;
cos[2613]=-6;
cos[2614]=-6;
cos[2615]=-6;
cos[2616]=-6;
cos[2617]=-6;
cos[2618]=-6;
cos[2619]=-6;
cos[2620]=-6;
cos[2621]=-6;
cos[2622]=-6;
cos[2623]=-6;
cos[2624]=-6;
cos[2625]=-6;
cos[2626]=-6;
cos[2627]=-6;
cos[2628]=-6;
cos[2629]=-6;
cos[2630]=-6;
cos[2631]=-6;
cos[2632]=-6;
cos[2633]=-7;
cos[2634]=-7;
cos[2635]=-7;
cos[2636]=-7;
cos[2637]=-7;
cos[2638]=-7;
cos[2639]=-7;
cos[2640]=-7;
cos[2641]=-7;
cos[2642]=-7;
cos[2643]=-7;
cos[2644]=-7;
cos[2645]=-7;
cos[2646]=-7;
cos[2647]=-7;
cos[2648]=-7;
cos[2649]=-7;
cos[2650]=-7;
cos[2651]=-7;
cos[2652]=-7;
cos[2653]=-7;
cos[2654]=-8;
cos[2655]=-8;
cos[2656]=-8;
cos[2657]=-8;
cos[2658]=-8;
cos[2659]=-8;
cos[2660]=-8;
cos[2661]=-8;
cos[2662]=-8;
cos[2663]=-8;
cos[2664]=-8;
cos[2665]=-8;
cos[2666]=-8;
cos[2667]=-8;
cos[2668]=-8;
cos[2669]=-8;
cos[2670]=-8;
cos[2671]=-8;
cos[2672]=-8;
cos[2673]=-8;
cos[2674]=-9;
cos[2675]=-9;
cos[2676]=-9;
cos[2677]=-9;
cos[2678]=-9;
cos[2679]=-9;
cos[2680]=-9;
cos[2681]=-9;
cos[2682]=-9;
cos[2683]=-9;
cos[2684]=-9;
cos[2685]=-9;
cos[2686]=-9;
cos[2687]=-9;
cos[2688]=-9;
cos[2689]=-9;
cos[2690]=-9;
cos[2691]=-9;
cos[2692]=-9;
cos[2693]=-9;
cos[2694]=-9;
cos[2695]=-10;
cos[2696]=-10;
cos[2697]=-10;
cos[2698]=-10;
cos[2699]=-10;
cos[2700]=-10;
cos[2701]=-10;
cos[2702]=-10;
cos[2703]=-10;
cos[2704]=-10;
cos[2705]=-10;
cos[2706]=-10;
cos[2707]=-10;
cos[2708]=-10;
cos[2709]=-10;
cos[2710]=-10;
cos[2711]=-10;
cos[2712]=-10;
cos[2713]=-10;
cos[2714]=-10;
cos[2715]=-11;
cos[2716]=-11;
cos[2717]=-11;
cos[2718]=-11;
cos[2719]=-11;
cos[2720]=-11;
cos[2721]=-11;
cos[2722]=-11;
cos[2723]=-11;
cos[2724]=-11;
cos[2725]=-11;
cos[2726]=-11;
cos[2727]=-11;
cos[2728]=-11;
cos[2729]=-11;
cos[2730]=-11;
cos[2731]=-11;
cos[2732]=-11;
cos[2733]=-11;
cos[2734]=-11;
cos[2735]=-11;
cos[2736]=-12;
cos[2737]=-12;
cos[2738]=-12;
cos[2739]=-12;
cos[2740]=-12;
cos[2741]=-12;
cos[2742]=-12;
cos[2743]=-12;
cos[2744]=-12;
cos[2745]=-12;
cos[2746]=-12;
cos[2747]=-12;
cos[2748]=-12;
cos[2749]=-12;
cos[2750]=-12;
cos[2751]=-12;
cos[2752]=-12;
cos[2753]=-12;
cos[2754]=-12;
cos[2755]=-12;
cos[2756]=-13;
cos[2757]=-13;
cos[2758]=-13;
cos[2759]=-13;
cos[2760]=-13;
cos[2761]=-13;
cos[2762]=-13;
cos[2763]=-13;
cos[2764]=-13;
cos[2765]=-13;
cos[2766]=-13;
cos[2767]=-13;
cos[2768]=-13;
cos[2769]=-13;
cos[2770]=-13;
cos[2771]=-13;
cos[2772]=-13;
cos[2773]=-13;
cos[2774]=-13;
cos[2775]=-13;
cos[2776]=-13;
cos[2777]=-14;
cos[2778]=-14;
cos[2779]=-14;
cos[2780]=-14;
cos[2781]=-14;
cos[2782]=-14;
cos[2783]=-14;
cos[2784]=-14;
cos[2785]=-14;
cos[2786]=-14;
cos[2787]=-14;
cos[2788]=-14;
cos[2789]=-14;
cos[2790]=-14;
cos[2791]=-14;
cos[2792]=-14;
cos[2793]=-14;
cos[2794]=-14;
cos[2795]=-14;
cos[2796]=-14;
cos[2797]=-14;
cos[2798]=-15;
cos[2799]=-15;
cos[2800]=-15;
cos[2801]=-15;
cos[2802]=-15;
cos[2803]=-15;
cos[2804]=-15;
cos[2805]=-15;
cos[2806]=-15;
cos[2807]=-15;
cos[2808]=-15;
cos[2809]=-15;
cos[2810]=-15;
cos[2811]=-15;
cos[2812]=-15;
cos[2813]=-15;
cos[2814]=-15;
cos[2815]=-15;
cos[2816]=-15;
cos[2817]=-15;
cos[2818]=-16;
cos[2819]=-16;
cos[2820]=-16;
cos[2821]=-16;
cos[2822]=-16;
cos[2823]=-16;
cos[2824]=-16;
cos[2825]=-16;
cos[2826]=-16;
cos[2827]=-16;
cos[2828]=-16;
cos[2829]=-16;
cos[2830]=-16;
cos[2831]=-16;
cos[2832]=-16;
cos[2833]=-16;
cos[2834]=-16;
cos[2835]=-16;
cos[2836]=-16;
cos[2837]=-16;
cos[2838]=-16;
cos[2839]=-17;
cos[2840]=-17;
cos[2841]=-17;
cos[2842]=-17;
cos[2843]=-17;
cos[2844]=-17;
cos[2845]=-17;
cos[2846]=-17;
cos[2847]=-17;
cos[2848]=-17;
cos[2849]=-17;
cos[2850]=-17;
cos[2851]=-17;
cos[2852]=-17;
cos[2853]=-17;
cos[2854]=-17;
cos[2855]=-17;
cos[2856]=-17;
cos[2857]=-17;
cos[2858]=-17;
cos[2859]=-17;
cos[2860]=-18;
cos[2861]=-18;
cos[2862]=-18;
cos[2863]=-18;
cos[2864]=-18;
cos[2865]=-18;
cos[2866]=-18;
cos[2867]=-18;
cos[2868]=-18;
cos[2869]=-18;
cos[2870]=-18;
cos[2871]=-18;
cos[2872]=-18;
cos[2873]=-18;
cos[2874]=-18;
cos[2875]=-18;
cos[2876]=-18;
cos[2877]=-18;
cos[2878]=-18;
cos[2879]=-18;
cos[2880]=-18;
cos[2881]=-19;
cos[2882]=-19;
cos[2883]=-19;
cos[2884]=-19;
cos[2885]=-19;
cos[2886]=-19;
cos[2887]=-19;
cos[2888]=-19;
cos[2889]=-19;
cos[2890]=-19;
cos[2891]=-19;
cos[2892]=-19;
cos[2893]=-19;
cos[2894]=-19;
cos[2895]=-19;
cos[2896]=-19;
cos[2897]=-19;
cos[2898]=-19;
cos[2899]=-19;
cos[2900]=-19;
cos[2901]=-19;
cos[2902]=-20;
cos[2903]=-20;
cos[2904]=-20;
cos[2905]=-20;
cos[2906]=-20;
cos[2907]=-20;
cos[2908]=-20;
cos[2909]=-20;
cos[2910]=-20;
cos[2911]=-20;
cos[2912]=-20;
cos[2913]=-20;
cos[2914]=-20;
cos[2915]=-20;
cos[2916]=-20;
cos[2917]=-20;
cos[2918]=-20;
cos[2919]=-20;
cos[2920]=-20;
cos[2921]=-20;
cos[2922]=-20;
cos[2923]=-21;
cos[2924]=-21;
cos[2925]=-21;
cos[2926]=-21;
cos[2927]=-21;
cos[2928]=-21;
cos[2929]=-21;
cos[2930]=-21;
cos[2931]=-21;
cos[2932]=-21;
cos[2933]=-21;
cos[2934]=-21;
cos[2935]=-21;
cos[2936]=-21;
cos[2937]=-21;
cos[2938]=-21;
cos[2939]=-21;
cos[2940]=-21;
cos[2941]=-21;
cos[2942]=-21;
cos[2943]=-21;
cos[2944]=-22;
cos[2945]=-22;
cos[2946]=-22;
cos[2947]=-22;
cos[2948]=-22;
cos[2949]=-22;
cos[2950]=-22;
cos[2951]=-22;
cos[2952]=-22;
cos[2953]=-22;
cos[2954]=-22;
cos[2955]=-22;
cos[2956]=-22;
cos[2957]=-22;
cos[2958]=-22;
cos[2959]=-22;
cos[2960]=-22;
cos[2961]=-22;
cos[2962]=-22;
cos[2963]=-22;
cos[2964]=-22;
cos[2965]=-23;
cos[2966]=-23;
cos[2967]=-23;
cos[2968]=-23;
cos[2969]=-23;
cos[2970]=-23;
cos[2971]=-23;
cos[2972]=-23;
cos[2973]=-23;
cos[2974]=-23;
cos[2975]=-23;
cos[2976]=-23;
cos[2977]=-23;
cos[2978]=-23;
cos[2979]=-23;
cos[2980]=-23;
cos[2981]=-23;
cos[2982]=-23;
cos[2983]=-23;
cos[2984]=-23;
cos[2985]=-23;
cos[2986]=-23;
cos[2987]=-24;
cos[2988]=-24;
cos[2989]=-24;
cos[2990]=-24;
cos[2991]=-24;
cos[2992]=-24;
cos[2993]=-24;
cos[2994]=-24;
cos[2995]=-24;
cos[2996]=-24;
cos[2997]=-24;
cos[2998]=-24;
cos[2999]=-24;
cos[3000]=-24;
cos[3001]=-24;
cos[3002]=-24;
cos[3003]=-24;
cos[3004]=-24;
cos[3005]=-24;
cos[3006]=-24;
cos[3007]=-24;
cos[3008]=-25;
cos[3009]=-25;
cos[3010]=-25;
cos[3011]=-25;
cos[3012]=-25;
cos[3013]=-25;
cos[3014]=-25;
cos[3015]=-25;
cos[3016]=-25;
cos[3017]=-25;
cos[3018]=-25;
cos[3019]=-25;
cos[3020]=-25;
cos[3021]=-25;
cos[3022]=-25;
cos[3023]=-25;
cos[3024]=-25;
cos[3025]=-25;
cos[3026]=-25;
cos[3027]=-25;
cos[3028]=-25;
cos[3029]=-25;
cos[3030]=-26;
cos[3031]=-26;
cos[3032]=-26;
cos[3033]=-26;
cos[3034]=-26;
cos[3035]=-26;
cos[3036]=-26;
cos[3037]=-26;
cos[3038]=-26;
cos[3039]=-26;
cos[3040]=-26;
cos[3041]=-26;
cos[3042]=-26;
cos[3043]=-26;
cos[3044]=-26;
cos[3045]=-26;
cos[3046]=-26;
cos[3047]=-26;
cos[3048]=-26;
cos[3049]=-26;
cos[3050]=-26;
cos[3051]=-27;
cos[3052]=-27;
cos[3053]=-27;
cos[3054]=-27;
cos[3055]=-27;
cos[3056]=-27;
cos[3057]=-27;
cos[3058]=-27;
cos[3059]=-27;
cos[3060]=-27;
cos[3061]=-27;
cos[3062]=-27;
cos[3063]=-27;
cos[3064]=-27;
cos[3065]=-27;
cos[3066]=-27;
cos[3067]=-27;
cos[3068]=-27;
cos[3069]=-27;
cos[3070]=-27;
cos[3071]=-27;
cos[3072]=-27;
cos[3073]=-28;
cos[3074]=-28;
cos[3075]=-28;
cos[3076]=-28;
cos[3077]=-28;
cos[3078]=-28;
cos[3079]=-28;
cos[3080]=-28;
cos[3081]=-28;
cos[3082]=-28;
cos[3083]=-28;
cos[3084]=-28;
cos[3085]=-28;
cos[3086]=-28;
cos[3087]=-28;
cos[3088]=-28;
cos[3089]=-28;
cos[3090]=-28;
cos[3091]=-28;
cos[3092]=-28;
cos[3093]=-28;
cos[3094]=-28;
cos[3095]=-29;
cos[3096]=-29;
cos[3097]=-29;
cos[3098]=-29;
cos[3099]=-29;
cos[3100]=-29;
cos[3101]=-29;
cos[3102]=-29;
cos[3103]=-29;
cos[3104]=-29;
cos[3105]=-29;
cos[3106]=-29;
cos[3107]=-29;
cos[3108]=-29;
cos[3109]=-29;
cos[3110]=-29;
cos[3111]=-29;
cos[3112]=-29;
cos[3113]=-29;
cos[3114]=-29;
cos[3115]=-29;
cos[3116]=-29;
cos[3117]=-30;
cos[3118]=-30;
cos[3119]=-30;
cos[3120]=-30;
cos[3121]=-30;
cos[3122]=-30;
cos[3123]=-30;
cos[3124]=-30;
cos[3125]=-30;
cos[3126]=-30;
cos[3127]=-30;
cos[3128]=-30;
cos[3129]=-30;
cos[3130]=-30;
cos[3131]=-30;
cos[3132]=-30;
cos[3133]=-30;
cos[3134]=-30;
cos[3135]=-30;
cos[3136]=-30;
cos[3137]=-30;
cos[3138]=-30;
cos[3139]=-31;
cos[3140]=-31;
cos[3141]=-31;
cos[3142]=-31;
cos[3143]=-31;
cos[3144]=-31;
cos[3145]=-31;
cos[3146]=-31;
cos[3147]=-31;
cos[3148]=-31;
cos[3149]=-31;
cos[3150]=-31;
cos[3151]=-31;
cos[3152]=-31;
cos[3153]=-31;
cos[3154]=-31;
cos[3155]=-31;
cos[3156]=-31;
cos[3157]=-31;
cos[3158]=-31;
cos[3159]=-31;
cos[3160]=-31;
cos[3161]=-32;
cos[3162]=-32;
cos[3163]=-32;
cos[3164]=-32;
cos[3165]=-32;
cos[3166]=-32;
cos[3167]=-32;
cos[3168]=-32;
cos[3169]=-32;
cos[3170]=-32;
cos[3171]=-32;
cos[3172]=-32;
cos[3173]=-32;
cos[3174]=-32;
cos[3175]=-32;
cos[3176]=-32;
cos[3177]=-32;
cos[3178]=-32;
cos[3179]=-32;
cos[3180]=-32;
cos[3181]=-32;
cos[3182]=-32;
cos[3183]=-33;
cos[3184]=-33;
cos[3185]=-33;
cos[3186]=-33;
cos[3187]=-33;
cos[3188]=-33;
cos[3189]=-33;
cos[3190]=-33;
cos[3191]=-33;
cos[3192]=-33;
cos[3193]=-33;
cos[3194]=-33;
cos[3195]=-33;
cos[3196]=-33;
cos[3197]=-33;
cos[3198]=-33;
cos[3199]=-33;
cos[3200]=-33;
cos[3201]=-33;
cos[3202]=-33;
cos[3203]=-33;
cos[3204]=-33;
cos[3205]=-33;
cos[3206]=-34;
cos[3207]=-34;
cos[3208]=-34;
cos[3209]=-34;
cos[3210]=-34;
cos[3211]=-34;
cos[3212]=-34;
cos[3213]=-34;
cos[3214]=-34;
cos[3215]=-34;
cos[3216]=-34;
cos[3217]=-34;
cos[3218]=-34;
cos[3219]=-34;
cos[3220]=-34;
cos[3221]=-34;
cos[3222]=-34;
cos[3223]=-34;
cos[3224]=-34;
cos[3225]=-34;
cos[3226]=-34;
cos[3227]=-34;
cos[3228]=-35;
cos[3229]=-35;
cos[3230]=-35;
cos[3231]=-35;
cos[3232]=-35;
cos[3233]=-35;
cos[3234]=-35;
cos[3235]=-35;
cos[3236]=-35;
cos[3237]=-35;
cos[3238]=-35;
cos[3239]=-35;
cos[3240]=-35;
cos[3241]=-35;
cos[3242]=-35;
cos[3243]=-35;
cos[3244]=-35;
cos[3245]=-35;
cos[3246]=-35;
cos[3247]=-35;
cos[3248]=-35;
cos[3249]=-35;
cos[3250]=-35;
cos[3251]=-36;
cos[3252]=-36;
cos[3253]=-36;
cos[3254]=-36;
cos[3255]=-36;
cos[3256]=-36;
cos[3257]=-36;
cos[3258]=-36;
cos[3259]=-36;
cos[3260]=-36;
cos[3261]=-36;
cos[3262]=-36;
cos[3263]=-36;
cos[3264]=-36;
cos[3265]=-36;
cos[3266]=-36;
cos[3267]=-36;
cos[3268]=-36;
cos[3269]=-36;
cos[3270]=-36;
cos[3271]=-36;
cos[3272]=-36;
cos[3273]=-36;
cos[3274]=-37;
cos[3275]=-37;
cos[3276]=-37;
cos[3277]=-37;
cos[3278]=-37;
cos[3279]=-37;
cos[3280]=-37;
cos[3281]=-37;
cos[3282]=-37;
cos[3283]=-37;
cos[3284]=-37;
cos[3285]=-37;
cos[3286]=-37;
cos[3287]=-37;
cos[3288]=-37;
cos[3289]=-37;
cos[3290]=-37;
cos[3291]=-37;
cos[3292]=-37;
cos[3293]=-37;
cos[3294]=-37;
cos[3295]=-37;
cos[3296]=-37;
cos[3297]=-38;
cos[3298]=-38;
cos[3299]=-38;
cos[3300]=-38;
cos[3301]=-38;
cos[3302]=-38;
cos[3303]=-38;
cos[3304]=-38;
cos[3305]=-38;
cos[3306]=-38;
cos[3307]=-38;
cos[3308]=-38;
cos[3309]=-38;
cos[3310]=-38;
cos[3311]=-38;
cos[3312]=-38;
cos[3313]=-38;
cos[3314]=-38;
cos[3315]=-38;
cos[3316]=-38;
cos[3317]=-38;
cos[3318]=-38;
cos[3319]=-38;
cos[3320]=-38;
cos[3321]=-39;
cos[3322]=-39;
cos[3323]=-39;
cos[3324]=-39;
cos[3325]=-39;
cos[3326]=-39;
cos[3327]=-39;
cos[3328]=-39;
cos[3329]=-39;
cos[3330]=-39;
cos[3331]=-39;
cos[3332]=-39;
cos[3333]=-39;
cos[3334]=-39;
cos[3335]=-39;
cos[3336]=-39;
cos[3337]=-39;
cos[3338]=-39;
cos[3339]=-39;
cos[3340]=-39;
cos[3341]=-39;
cos[3342]=-39;
cos[3343]=-39;
cos[3344]=-40;
cos[3345]=-40;
cos[3346]=-40;
cos[3347]=-40;
cos[3348]=-40;
cos[3349]=-40;
cos[3350]=-40;
cos[3351]=-40;
cos[3352]=-40;
cos[3353]=-40;
cos[3354]=-40;
cos[3355]=-40;
cos[3356]=-40;
cos[3357]=-40;
cos[3358]=-40;
cos[3359]=-40;
cos[3360]=-40;
cos[3361]=-40;
cos[3362]=-40;
cos[3363]=-40;
cos[3364]=-40;
cos[3365]=-40;
cos[3366]=-40;
cos[3367]=-40;
cos[3368]=-41;
cos[3369]=-41;
cos[3370]=-41;
cos[3371]=-41;
cos[3372]=-41;
cos[3373]=-41;
cos[3374]=-41;
cos[3375]=-41;
cos[3376]=-41;
cos[3377]=-41;
cos[3378]=-41;
cos[3379]=-41;
cos[3380]=-41;
cos[3381]=-41;
cos[3382]=-41;
cos[3383]=-41;
cos[3384]=-41;
cos[3385]=-41;
cos[3386]=-41;
cos[3387]=-41;
cos[3388]=-41;
cos[3389]=-41;
cos[3390]=-41;
cos[3391]=-41;
cos[3392]=-42;
cos[3393]=-42;
cos[3394]=-42;
cos[3395]=-42;
cos[3396]=-42;
cos[3397]=-42;
cos[3398]=-42;
cos[3399]=-42;
cos[3400]=-42;
cos[3401]=-42;
cos[3402]=-42;
cos[3403]=-42;
cos[3404]=-42;
cos[3405]=-42;
cos[3406]=-42;
cos[3407]=-42;
cos[3408]=-42;
cos[3409]=-42;
cos[3410]=-42;
cos[3411]=-42;
cos[3412]=-42;
cos[3413]=-42;
cos[3414]=-42;
cos[3415]=-42;
cos[3416]=-43;
cos[3417]=-43;
cos[3418]=-43;
cos[3419]=-43;
cos[3420]=-43;
cos[3421]=-43;
cos[3422]=-43;
cos[3423]=-43;
cos[3424]=-43;
cos[3425]=-43;
cos[3426]=-43;
cos[3427]=-43;
cos[3428]=-43;
cos[3429]=-43;
cos[3430]=-43;
cos[3431]=-43;
cos[3432]=-43;
cos[3433]=-43;
cos[3434]=-43;
cos[3435]=-43;
cos[3436]=-43;
cos[3437]=-43;
cos[3438]=-43;
cos[3439]=-43;
cos[3440]=-44;
cos[3441]=-44;
cos[3442]=-44;
cos[3443]=-44;
cos[3444]=-44;
cos[3445]=-44;
cos[3446]=-44;
cos[3447]=-44;
cos[3448]=-44;
cos[3449]=-44;
cos[3450]=-44;
cos[3451]=-44;
cos[3452]=-44;
cos[3453]=-44;
cos[3454]=-44;
cos[3455]=-44;
cos[3456]=-44;
cos[3457]=-44;
cos[3458]=-44;
cos[3459]=-44;
cos[3460]=-44;
cos[3461]=-44;
cos[3462]=-44;
cos[3463]=-44;
cos[3464]=-44;
cos[3465]=-45;
cos[3466]=-45;
cos[3467]=-45;
cos[3468]=-45;
cos[3469]=-45;
cos[3470]=-45;
cos[3471]=-45;
cos[3472]=-45;
cos[3473]=-45;
cos[3474]=-45;
cos[3475]=-45;
cos[3476]=-45;
cos[3477]=-45;
cos[3478]=-45;
cos[3479]=-45;
cos[3480]=-45;
cos[3481]=-45;
cos[3482]=-45;
cos[3483]=-45;
cos[3484]=-45;
cos[3485]=-45;
cos[3486]=-45;
cos[3487]=-45;
cos[3488]=-45;
cos[3489]=-45;
cos[3490]=-46;
cos[3491]=-46;
cos[3492]=-46;
cos[3493]=-46;
cos[3494]=-46;
cos[3495]=-46;
cos[3496]=-46;
cos[3497]=-46;
cos[3498]=-46;
cos[3499]=-46;
cos[3500]=-46;
cos[3501]=-46;
cos[3502]=-46;
cos[3503]=-46;
cos[3504]=-46;
cos[3505]=-46;
cos[3506]=-46;
cos[3507]=-46;
cos[3508]=-46;
cos[3509]=-46;
cos[3510]=-46;
cos[3511]=-46;
cos[3512]=-46;
cos[3513]=-46;
cos[3514]=-46;
cos[3515]=-47;
cos[3516]=-47;
cos[3517]=-47;
cos[3518]=-47;
cos[3519]=-47;
cos[3520]=-47;
cos[3521]=-47;
cos[3522]=-47;
cos[3523]=-47;
cos[3524]=-47;
cos[3525]=-47;
cos[3526]=-47;
cos[3527]=-47;
cos[3528]=-47;
cos[3529]=-47;
cos[3530]=-47;
cos[3531]=-47;
cos[3532]=-47;
cos[3533]=-47;
cos[3534]=-47;
cos[3535]=-47;
cos[3536]=-47;
cos[3537]=-47;
cos[3538]=-47;
cos[3539]=-47;
cos[3540]=-47;
cos[3541]=-48;
cos[3542]=-48;
cos[3543]=-48;
cos[3544]=-48;
cos[3545]=-48;
cos[3546]=-48;
cos[3547]=-48;
cos[3548]=-48;
cos[3549]=-48;
cos[3550]=-48;
cos[3551]=-48;
cos[3552]=-48;
cos[3553]=-48;
cos[3554]=-48;
cos[3555]=-48;
cos[3556]=-48;
cos[3557]=-48;
cos[3558]=-48;
cos[3559]=-48;
cos[3560]=-48;
cos[3561]=-48;
cos[3562]=-48;
cos[3563]=-48;
cos[3564]=-48;
cos[3565]=-48;
cos[3566]=-49;
cos[3567]=-49;
cos[3568]=-49;
cos[3569]=-49;
cos[3570]=-49;
cos[3571]=-49;
cos[3572]=-49;
cos[3573]=-49;
cos[3574]=-49;
cos[3575]=-49;
cos[3576]=-49;
cos[3577]=-49;
cos[3578]=-49;
cos[3579]=-49;
cos[3580]=-49;
cos[3581]=-49;
cos[3582]=-49;
cos[3583]=-49;
cos[3584]=-49;
cos[3585]=-49;
cos[3586]=-49;
cos[3587]=-49;
cos[3588]=-49;
cos[3589]=-49;
cos[3590]=-49;
cos[3591]=-49;
cos[3592]=-49;
cos[3593]=-50;
cos[3594]=-50;
cos[3595]=-50;
cos[3596]=-50;
cos[3597]=-50;
cos[3598]=-50;
cos[3599]=-50;
cos[3600]=-50;
cos[3601]=-50;
cos[3602]=-50;
cos[3603]=-50;
cos[3604]=-50;
cos[3605]=-50;
cos[3606]=-50;
cos[3607]=-50;
cos[3608]=-50;
cos[3609]=-50;
cos[3610]=-50;
cos[3611]=-50;
cos[3612]=-50;
cos[3613]=-50;
cos[3614]=-50;
cos[3615]=-50;
cos[3616]=-50;
cos[3617]=-50;
cos[3618]=-50;
cos[3619]=-51;
cos[3620]=-51;
cos[3621]=-51;
cos[3622]=-51;
cos[3623]=-51;
cos[3624]=-51;
cos[3625]=-51;
cos[3626]=-51;
cos[3627]=-51;
cos[3628]=-51;
cos[3629]=-51;
cos[3630]=-51;
cos[3631]=-51;
cos[3632]=-51;
cos[3633]=-51;
cos[3634]=-51;
cos[3635]=-51;
cos[3636]=-51;
cos[3637]=-51;
cos[3638]=-51;
cos[3639]=-51;
cos[3640]=-51;
cos[3641]=-51;
cos[3642]=-51;
cos[3643]=-51;
cos[3644]=-51;
cos[3645]=-51;
cos[3646]=-52;
cos[3647]=-52;
cos[3648]=-52;
cos[3649]=-52;
cos[3650]=-52;
cos[3651]=-52;
cos[3652]=-52;
cos[3653]=-52;
cos[3654]=-52;
cos[3655]=-52;
cos[3656]=-52;
cos[3657]=-52;
cos[3658]=-52;
cos[3659]=-52;
cos[3660]=-52;
cos[3661]=-52;
cos[3662]=-52;
cos[3663]=-52;
cos[3664]=-52;
cos[3665]=-52;
cos[3666]=-52;
cos[3667]=-52;
cos[3668]=-52;
cos[3669]=-52;
cos[3670]=-52;
cos[3671]=-52;
cos[3672]=-52;
cos[3673]=-53;
cos[3674]=-53;
cos[3675]=-53;
cos[3676]=-53;
cos[3677]=-53;
cos[3678]=-53;
cos[3679]=-53;
cos[3680]=-53;
cos[3681]=-53;
cos[3682]=-53;
cos[3683]=-53;
cos[3684]=-53;
cos[3685]=-53;
cos[3686]=-53;
cos[3687]=-53;
cos[3688]=-53;
cos[3689]=-53;
cos[3690]=-53;
cos[3691]=-53;
cos[3692]=-53;
cos[3693]=-53;
cos[3694]=-53;
cos[3695]=-53;
cos[3696]=-53;
cos[3697]=-53;
cos[3698]=-53;
cos[3699]=-53;
cos[3700]=-53;
cos[3701]=-54;
cos[3702]=-54;
cos[3703]=-54;
cos[3704]=-54;
cos[3705]=-54;
cos[3706]=-54;
cos[3707]=-54;
cos[3708]=-54;
cos[3709]=-54;
cos[3710]=-54;
cos[3711]=-54;
cos[3712]=-54;
cos[3713]=-54;
cos[3714]=-54;
cos[3715]=-54;
cos[3716]=-54;
cos[3717]=-54;
cos[3718]=-54;
cos[3719]=-54;
cos[3720]=-54;
cos[3721]=-54;
cos[3722]=-54;
cos[3723]=-54;
cos[3724]=-54;
cos[3725]=-54;
cos[3726]=-54;
cos[3727]=-54;
cos[3728]=-54;
cos[3729]=-55;
cos[3730]=-55;
cos[3731]=-55;
cos[3732]=-55;
cos[3733]=-55;
cos[3734]=-55;
cos[3735]=-55;
cos[3736]=-55;
cos[3737]=-55;
cos[3738]=-55;
cos[3739]=-55;
cos[3740]=-55;
cos[3741]=-55;
cos[3742]=-55;
cos[3743]=-55;
cos[3744]=-55;
cos[3745]=-55;
cos[3746]=-55;
cos[3747]=-55;
cos[3748]=-55;
cos[3749]=-55;
cos[3750]=-55;
cos[3751]=-55;
cos[3752]=-55;
cos[3753]=-55;
cos[3754]=-55;
cos[3755]=-55;
cos[3756]=-55;
cos[3757]=-55;
cos[3758]=-56;
cos[3759]=-56;
cos[3760]=-56;
cos[3761]=-56;
cos[3762]=-56;
cos[3763]=-56;
cos[3764]=-56;
cos[3765]=-56;
cos[3766]=-56;
cos[3767]=-56;
cos[3768]=-56;
cos[3769]=-56;
cos[3770]=-56;
cos[3771]=-56;
cos[3772]=-56;
cos[3773]=-56;
cos[3774]=-56;
cos[3775]=-56;
cos[3776]=-56;
cos[3777]=-56;
cos[3778]=-56;
cos[3779]=-56;
cos[3780]=-56;
cos[3781]=-56;
cos[3782]=-56;
cos[3783]=-56;
cos[3784]=-56;
cos[3785]=-56;
cos[3786]=-56;
cos[3787]=-57;
cos[3788]=-57;
cos[3789]=-57;
cos[3790]=-57;
cos[3791]=-57;
cos[3792]=-57;
cos[3793]=-57;
cos[3794]=-57;
cos[3795]=-57;
cos[3796]=-57;
cos[3797]=-57;
cos[3798]=-57;
cos[3799]=-57;
cos[3800]=-57;
cos[3801]=-57;
cos[3802]=-57;
cos[3803]=-57;
cos[3804]=-57;
cos[3805]=-57;
cos[3806]=-57;
cos[3807]=-57;
cos[3808]=-57;
cos[3809]=-57;
cos[3810]=-57;
cos[3811]=-57;
cos[3812]=-57;
cos[3813]=-57;
cos[3814]=-57;
cos[3815]=-57;
cos[3816]=-57;
cos[3817]=-58;
cos[3818]=-58;
cos[3819]=-58;
cos[3820]=-58;
cos[3821]=-58;
cos[3822]=-58;
cos[3823]=-58;
cos[3824]=-58;
cos[3825]=-58;
cos[3826]=-58;
cos[3827]=-58;
cos[3828]=-58;
cos[3829]=-58;
cos[3830]=-58;
cos[3831]=-58;
cos[3832]=-58;
cos[3833]=-58;
cos[3834]=-58;
cos[3835]=-58;
cos[3836]=-58;
cos[3837]=-58;
cos[3838]=-58;
cos[3839]=-58;
cos[3840]=-58;
cos[3841]=-58;
cos[3842]=-58;
cos[3843]=-58;
cos[3844]=-58;
cos[3845]=-58;
cos[3846]=-58;
cos[3847]=-59;
cos[3848]=-59;
cos[3849]=-59;
cos[3850]=-59;
cos[3851]=-59;
cos[3852]=-59;
cos[3853]=-59;
cos[3854]=-59;
cos[3855]=-59;
cos[3856]=-59;
cos[3857]=-59;
cos[3858]=-59;
cos[3859]=-59;
cos[3860]=-59;
cos[3861]=-59;
cos[3862]=-59;
cos[3863]=-59;
cos[3864]=-59;
cos[3865]=-59;
cos[3866]=-59;
cos[3867]=-59;
cos[3868]=-59;
cos[3869]=-59;
cos[3870]=-59;
cos[3871]=-59;
cos[3872]=-59;
cos[3873]=-59;
cos[3874]=-59;
cos[3875]=-59;
cos[3876]=-59;
cos[3877]=-59;
cos[3878]=-60;
cos[3879]=-60;
cos[3880]=-60;
cos[3881]=-60;
cos[3882]=-60;
cos[3883]=-60;
cos[3884]=-60;
cos[3885]=-60;
cos[3886]=-60;
cos[3887]=-60;
cos[3888]=-60;
cos[3889]=-60;
cos[3890]=-60;
cos[3891]=-60;
cos[3892]=-60;
cos[3893]=-60;
cos[3894]=-60;
cos[3895]=-60;
cos[3896]=-60;
cos[3897]=-60;
cos[3898]=-60;
cos[3899]=-60;
cos[3900]=-60;
cos[3901]=-60;
cos[3902]=-60;
cos[3903]=-60;
cos[3904]=-60;
cos[3905]=-60;
cos[3906]=-60;
cos[3907]=-60;
cos[3908]=-60;
cos[3909]=-60;
cos[3910]=-61;
cos[3911]=-61;
cos[3912]=-61;
cos[3913]=-61;
cos[3914]=-61;
cos[3915]=-61;
cos[3916]=-61;
cos[3917]=-61;
cos[3918]=-61;
cos[3919]=-61;
cos[3920]=-61;
cos[3921]=-61;
cos[3922]=-61;
cos[3923]=-61;
cos[3924]=-61;
cos[3925]=-61;
cos[3926]=-61;
cos[3927]=-61;
cos[3928]=-61;
cos[3929]=-61;
cos[3930]=-61;
cos[3931]=-61;
cos[3932]=-61;
cos[3933]=-61;
cos[3934]=-61;
cos[3935]=-61;
cos[3936]=-61;
cos[3937]=-61;
cos[3938]=-61;
cos[3939]=-61;
cos[3940]=-61;
cos[3941]=-61;
cos[3942]=-61;
cos[3943]=-62;
cos[3944]=-62;
cos[3945]=-62;
cos[3946]=-62;
cos[3947]=-62;
cos[3948]=-62;
cos[3949]=-62;
cos[3950]=-62;
cos[3951]=-62;
cos[3952]=-62;
cos[3953]=-62;
cos[3954]=-62;
cos[3955]=-62;
cos[3956]=-62;
cos[3957]=-62;
cos[3958]=-62;
cos[3959]=-62;
cos[3960]=-62;
cos[3961]=-62;
cos[3962]=-62;
cos[3963]=-62;
cos[3964]=-62;
cos[3965]=-62;
cos[3966]=-62;
cos[3967]=-62;
cos[3968]=-62;
cos[3969]=-62;
cos[3970]=-62;
cos[3971]=-62;
cos[3972]=-62;
cos[3973]=-62;
cos[3974]=-62;
cos[3975]=-62;
cos[3976]=-63;
cos[3977]=-63;
cos[3978]=-63;
cos[3979]=-63;
cos[3980]=-63;
cos[3981]=-63;
cos[3982]=-63;
cos[3983]=-63;
cos[3984]=-63;
cos[3985]=-63;
cos[3986]=-63;
cos[3987]=-63;
cos[3988]=-63;
cos[3989]=-63;
cos[3990]=-63;
cos[3991]=-63;
cos[3992]=-63;
cos[3993]=-63;
cos[3994]=-63;
cos[3995]=-63;
cos[3996]=-63;
cos[3997]=-63;
cos[3998]=-63;
cos[3999]=-63;
cos[4000]=-63;
cos[4001]=-63;
cos[4002]=-63;
cos[4003]=-63;
cos[4004]=-63;
cos[4005]=-63;
cos[4006]=-63;
cos[4007]=-63;
cos[4008]=-63;
cos[4009]=-63;
cos[4010]=-63;
cos[4011]=-64;
cos[4012]=-64;
cos[4013]=-64;
cos[4014]=-64;
cos[4015]=-64;
cos[4016]=-64;
cos[4017]=-64;
cos[4018]=-64;
cos[4019]=-64;
cos[4020]=-64;
cos[4021]=-64;
cos[4022]=-64;
cos[4023]=-64;
cos[4024]=-64;
cos[4025]=-64;
cos[4026]=-64;
cos[4027]=-64;
cos[4028]=-64;
cos[4029]=-64;
cos[4030]=-64;
cos[4031]=-64;
cos[4032]=-64;
cos[4033]=-64;
cos[4034]=-64;
cos[4035]=-64;
cos[4036]=-64;
cos[4037]=-64;
cos[4038]=-64;
cos[4039]=-64;
cos[4040]=-64;
cos[4041]=-64;
cos[4042]=-64;
cos[4043]=-64;
cos[4044]=-64;
cos[4045]=-64;
cos[4046]=-65;
cos[4047]=-65;
cos[4048]=-65;
cos[4049]=-65;
cos[4050]=-65;
cos[4051]=-65;
cos[4052]=-65;
cos[4053]=-65;
cos[4054]=-65;
cos[4055]=-65;
cos[4056]=-65;
cos[4057]=-65;
cos[4058]=-65;
cos[4059]=-65;
cos[4060]=-65;
cos[4061]=-65;
cos[4062]=-65;
cos[4063]=-65;
cos[4064]=-65;
cos[4065]=-65;
cos[4066]=-65;
cos[4067]=-65;
cos[4068]=-65;
cos[4069]=-65;
cos[4070]=-65;
cos[4071]=-65;
cos[4072]=-65;
cos[4073]=-65;
cos[4074]=-65;
cos[4075]=-65;
cos[4076]=-65;
cos[4077]=-65;
cos[4078]=-65;
cos[4079]=-65;
cos[4080]=-65;
cos[4081]=-65;
cos[4082]=-65;
cos[4083]=-66;
cos[4084]=-66;
cos[4085]=-66;
cos[4086]=-66;
cos[4087]=-66;
cos[4088]=-66;
cos[4089]=-66;
cos[4090]=-66;
cos[4091]=-66;
cos[4092]=-66;
cos[4093]=-66;
cos[4094]=-66;
cos[4095]=-66;
cos[4096]=-66;
cos[4097]=-66;
cos[4098]=-66;
cos[4099]=-66;
cos[4100]=-66;
cos[4101]=-66;
cos[4102]=-66;
cos[4103]=-66;
cos[4104]=-66;
cos[4105]=-66;
cos[4106]=-66;
cos[4107]=-66;
cos[4108]=-66;
cos[4109]=-66;
cos[4110]=-66;
cos[4111]=-66;
cos[4112]=-66;
cos[4113]=-66;
cos[4114]=-66;
cos[4115]=-66;
cos[4116]=-66;
cos[4117]=-66;
cos[4118]=-66;
cos[4119]=-66;
cos[4120]=-66;
cos[4121]=-67;
cos[4122]=-67;
cos[4123]=-67;
cos[4124]=-67;
cos[4125]=-67;
cos[4126]=-67;
cos[4127]=-67;
cos[4128]=-67;
cos[4129]=-67;
cos[4130]=-67;
cos[4131]=-67;
cos[4132]=-67;
cos[4133]=-67;
cos[4134]=-67;
cos[4135]=-67;
cos[4136]=-67;
cos[4137]=-67;
cos[4138]=-67;
cos[4139]=-67;
cos[4140]=-67;
cos[4141]=-67;
cos[4142]=-67;
cos[4143]=-67;
cos[4144]=-67;
cos[4145]=-67;
cos[4146]=-67;
cos[4147]=-67;
cos[4148]=-67;
cos[4149]=-67;
cos[4150]=-67;
cos[4151]=-67;
cos[4152]=-67;
cos[4153]=-67;
cos[4154]=-67;
cos[4155]=-67;
cos[4156]=-67;
cos[4157]=-67;
cos[4158]=-67;
cos[4159]=-67;
cos[4160]=-67;
cos[4161]=-68;
cos[4162]=-68;
cos[4163]=-68;
cos[4164]=-68;
cos[4165]=-68;
cos[4166]=-68;
cos[4167]=-68;
cos[4168]=-68;
cos[4169]=-68;
cos[4170]=-68;
cos[4171]=-68;
cos[4172]=-68;
cos[4173]=-68;
cos[4174]=-68;
cos[4175]=-68;
cos[4176]=-68;
cos[4177]=-68;
cos[4178]=-68;
cos[4179]=-68;
cos[4180]=-68;
cos[4181]=-68;
cos[4182]=-68;
cos[4183]=-68;
cos[4184]=-68;
cos[4185]=-68;
cos[4186]=-68;
cos[4187]=-68;
cos[4188]=-68;
cos[4189]=-68;
cos[4190]=-68;
cos[4191]=-68;
cos[4192]=-68;
cos[4193]=-68;
cos[4194]=-68;
cos[4195]=-68;
cos[4196]=-68;
cos[4197]=-68;
cos[4198]=-68;
cos[4199]=-68;
cos[4200]=-68;
cos[4201]=-68;
cos[4202]=-69;
cos[4203]=-69;
cos[4204]=-69;
cos[4205]=-69;
cos[4206]=-69;
cos[4207]=-69;
cos[4208]=-69;
cos[4209]=-69;
cos[4210]=-69;
cos[4211]=-69;
cos[4212]=-69;
cos[4213]=-69;
cos[4214]=-69;
cos[4215]=-69;
cos[4216]=-69;
cos[4217]=-69;
cos[4218]=-69;
cos[4219]=-69;
cos[4220]=-69;
cos[4221]=-69;
cos[4222]=-69;
cos[4223]=-69;
cos[4224]=-69;
cos[4225]=-69;
cos[4226]=-69;
cos[4227]=-69;
cos[4228]=-69;
cos[4229]=-69;
cos[4230]=-69;
cos[4231]=-69;
cos[4232]=-69;
cos[4233]=-69;
cos[4234]=-69;
cos[4235]=-69;
cos[4236]=-69;
cos[4237]=-69;
cos[4238]=-69;
cos[4239]=-69;
cos[4240]=-69;
cos[4241]=-69;
cos[4242]=-69;
cos[4243]=-69;
cos[4244]=-69;
cos[4245]=-69;
cos[4246]=-70;
cos[4247]=-70;
cos[4248]=-70;
cos[4249]=-70;
cos[4250]=-70;
cos[4251]=-70;
cos[4252]=-70;
cos[4253]=-70;
cos[4254]=-70;
cos[4255]=-70;
cos[4256]=-70;
cos[4257]=-70;
cos[4258]=-70;
cos[4259]=-70;
cos[4260]=-70;
cos[4261]=-70;
cos[4262]=-70;
cos[4263]=-70;
cos[4264]=-70;
cos[4265]=-70;
cos[4266]=-70;
cos[4267]=-70;
cos[4268]=-70;
cos[4269]=-70;
cos[4270]=-70;
cos[4271]=-70;
cos[4272]=-70;
cos[4273]=-70;
cos[4274]=-70;
cos[4275]=-70;
cos[4276]=-70;
cos[4277]=-70;
cos[4278]=-70;
cos[4279]=-70;
cos[4280]=-70;
cos[4281]=-70;
cos[4282]=-70;
cos[4283]=-70;
cos[4284]=-70;
cos[4285]=-70;
cos[4286]=-70;
cos[4287]=-70;
cos[4288]=-70;
cos[4289]=-70;
cos[4290]=-70;
cos[4291]=-71;
cos[4292]=-71;
cos[4293]=-71;
cos[4294]=-71;
cos[4295]=-71;
cos[4296]=-71;
cos[4297]=-71;
cos[4298]=-71;
cos[4299]=-71;
cos[4300]=-71;
cos[4301]=-71;
cos[4302]=-71;
cos[4303]=-71;
cos[4304]=-71;
cos[4305]=-71;
cos[4306]=-71;
cos[4307]=-71;
cos[4308]=-71;
cos[4309]=-71;
cos[4310]=-71;
cos[4311]=-71;
cos[4312]=-71;
cos[4313]=-71;
cos[4314]=-71;
cos[4315]=-71;
cos[4316]=-71;
cos[4317]=-71;
cos[4318]=-71;
cos[4319]=-71;
cos[4320]=-71;
cos[4321]=-71;
cos[4322]=-71;
cos[4323]=-71;
cos[4324]=-71;
cos[4325]=-71;
cos[4326]=-71;
cos[4327]=-71;
cos[4328]=-71;
cos[4329]=-71;
cos[4330]=-71;
cos[4331]=-71;
cos[4332]=-71;
cos[4333]=-71;
cos[4334]=-71;
cos[4335]=-71;
cos[4336]=-71;
cos[4337]=-71;
cos[4338]=-71;
cos[4339]=-71;
cos[4340]=-72;
cos[4341]=-72;
cos[4342]=-72;
cos[4343]=-72;
cos[4344]=-72;
cos[4345]=-72;
cos[4346]=-72;
cos[4347]=-72;
cos[4348]=-72;
cos[4349]=-72;
cos[4350]=-72;
cos[4351]=-72;
cos[4352]=-72;
cos[4353]=-72;
cos[4354]=-72;
cos[4355]=-72;
cos[4356]=-72;
cos[4357]=-72;
cos[4358]=-72;
cos[4359]=-72;
cos[4360]=-72;
cos[4361]=-72;
cos[4362]=-72;
cos[4363]=-72;
cos[4364]=-72;
cos[4365]=-72;
cos[4366]=-72;
cos[4367]=-72;
cos[4368]=-72;
cos[4369]=-72;
cos[4370]=-72;
cos[4371]=-72;
cos[4372]=-72;
cos[4373]=-72;
cos[4374]=-72;
cos[4375]=-72;
cos[4376]=-72;
cos[4377]=-72;
cos[4378]=-72;
cos[4379]=-72;
cos[4380]=-72;
cos[4381]=-72;
cos[4382]=-72;
cos[4383]=-72;
cos[4384]=-72;
cos[4385]=-72;
cos[4386]=-72;
cos[4387]=-72;
cos[4388]=-72;
cos[4389]=-72;
cos[4390]=-72;
cos[4391]=-72;
cos[4392]=-72;
cos[4393]=-73;
cos[4394]=-73;
cos[4395]=-73;
cos[4396]=-73;
cos[4397]=-73;
cos[4398]=-73;
cos[4399]=-73;
cos[4400]=-73;
cos[4401]=-73;
cos[4402]=-73;
cos[4403]=-73;
cos[4404]=-73;
cos[4405]=-73;
cos[4406]=-73;
cos[4407]=-73;
cos[4408]=-73;
cos[4409]=-73;
cos[4410]=-73;
cos[4411]=-73;
cos[4412]=-73;
cos[4413]=-73;
cos[4414]=-73;
cos[4415]=-73;
cos[4416]=-73;
cos[4417]=-73;
cos[4418]=-73;
cos[4419]=-73;
cos[4420]=-73;
cos[4421]=-73;
cos[4422]=-73;
cos[4423]=-73;
cos[4424]=-73;
cos[4425]=-73;
cos[4426]=-73;
cos[4427]=-73;
cos[4428]=-73;
cos[4429]=-73;
cos[4430]=-73;
cos[4431]=-73;
cos[4432]=-73;
cos[4433]=-73;
cos[4434]=-73;
cos[4435]=-73;
cos[4436]=-73;
cos[4437]=-73;
cos[4438]=-73;
cos[4439]=-73;
cos[4440]=-73;
cos[4441]=-73;
cos[4442]=-73;
cos[4443]=-73;
cos[4444]=-73;
cos[4445]=-73;
cos[4446]=-73;
cos[4447]=-73;
cos[4448]=-73;
cos[4449]=-73;
cos[4450]=-74;
cos[4451]=-74;
cos[4452]=-74;
cos[4453]=-74;
cos[4454]=-74;
cos[4455]=-74;
cos[4456]=-74;
cos[4457]=-74;
cos[4458]=-74;
cos[4459]=-74;
cos[4460]=-74;
cos[4461]=-74;
cos[4462]=-74;
cos[4463]=-74;
cos[4464]=-74;
cos[4465]=-74;
cos[4466]=-74;
cos[4467]=-74;
cos[4468]=-74;
cos[4469]=-74;
cos[4470]=-74;
cos[4471]=-74;
cos[4472]=-74;
cos[4473]=-74;
cos[4474]=-74;
cos[4475]=-74;
cos[4476]=-74;
cos[4477]=-74;
cos[4478]=-74;
cos[4479]=-74;
cos[4480]=-74;
cos[4481]=-74;
cos[4482]=-74;
cos[4483]=-74;
cos[4484]=-74;
cos[4485]=-74;
cos[4486]=-74;
cos[4487]=-74;
cos[4488]=-74;
cos[4489]=-74;
cos[4490]=-74;
cos[4491]=-74;
cos[4492]=-74;
cos[4493]=-74;
cos[4494]=-74;
cos[4495]=-74;
cos[4496]=-74;
cos[4497]=-74;
cos[4498]=-74;
cos[4499]=-74;
cos[4500]=-74;
cos[4501]=-74;
cos[4502]=-74;
cos[4503]=-74;
cos[4504]=-74;
cos[4505]=-74;
cos[4506]=-74;
cos[4507]=-74;
cos[4508]=-74;
cos[4509]=-74;
cos[4510]=-74;
cos[4511]=-74;
cos[4512]=-74;
cos[4513]=-74;
cos[4514]=-75;
cos[4515]=-75;
cos[4516]=-75;
cos[4517]=-75;
cos[4518]=-75;
cos[4519]=-75;
cos[4520]=-75;
cos[4521]=-75;
cos[4522]=-75;
cos[4523]=-75;
cos[4524]=-75;
cos[4525]=-75;
cos[4526]=-75;
cos[4527]=-75;
cos[4528]=-75;
cos[4529]=-75;
cos[4530]=-75;
cos[4531]=-75;
cos[4532]=-75;
cos[4533]=-75;
cos[4534]=-75;
cos[4535]=-75;
cos[4536]=-75;
cos[4537]=-75;
cos[4538]=-75;
cos[4539]=-75;
cos[4540]=-75;
cos[4541]=-75;
cos[4542]=-75;
cos[4543]=-75;
cos[4544]=-75;
cos[4545]=-75;
cos[4546]=-75;
cos[4547]=-75;
cos[4548]=-75;
cos[4549]=-75;
cos[4550]=-75;
cos[4551]=-75;
cos[4552]=-75;
cos[4553]=-75;
cos[4554]=-75;
cos[4555]=-75;
cos[4556]=-75;
cos[4557]=-75;
cos[4558]=-75;
cos[4559]=-75;
cos[4560]=-75;
cos[4561]=-75;
cos[4562]=-75;
cos[4563]=-75;
cos[4564]=-75;
cos[4565]=-75;
cos[4566]=-75;
cos[4567]=-75;
cos[4568]=-75;
cos[4569]=-75;
cos[4570]=-75;
cos[4571]=-75;
cos[4572]=-75;
cos[4573]=-75;
cos[4574]=-75;
cos[4575]=-75;
cos[4576]=-75;
cos[4577]=-75;
cos[4578]=-75;
cos[4579]=-75;
cos[4580]=-75;
cos[4581]=-75;
cos[4582]=-75;
cos[4583]=-75;
cos[4584]=-75;
cos[4585]=-75;
cos[4586]=-75;
cos[4587]=-76;
cos[4588]=-76;
cos[4589]=-76;
cos[4590]=-76;
cos[4591]=-76;
cos[4592]=-76;
cos[4593]=-76;
cos[4594]=-76;
cos[4595]=-76;
cos[4596]=-76;
cos[4597]=-76;
cos[4598]=-76;
cos[4599]=-76;
cos[4600]=-76;
cos[4601]=-76;
cos[4602]=-76;
cos[4603]=-76;
cos[4604]=-76;
cos[4605]=-76;
cos[4606]=-76;
cos[4607]=-76;
cos[4608]=-76;
cos[4609]=-76;
cos[4610]=-76;
cos[4611]=-76;
cos[4612]=-76;
cos[4613]=-76;
cos[4614]=-76;
cos[4615]=-76;
cos[4616]=-76;
cos[4617]=-76;
cos[4618]=-76;
cos[4619]=-76;
cos[4620]=-76;
cos[4621]=-76;
cos[4622]=-76;
cos[4623]=-76;
cos[4624]=-76;
cos[4625]=-76;
cos[4626]=-76;
cos[4627]=-76;
cos[4628]=-76;
cos[4629]=-76;
cos[4630]=-76;
cos[4631]=-76;
cos[4632]=-76;
cos[4633]=-76;
cos[4634]=-76;
cos[4635]=-76;
cos[4636]=-76;
cos[4637]=-76;
cos[4638]=-76;
cos[4639]=-76;
cos[4640]=-76;
cos[4641]=-76;
cos[4642]=-76;
cos[4643]=-76;
cos[4644]=-76;
cos[4645]=-76;
cos[4646]=-76;
cos[4647]=-76;
cos[4648]=-76;
cos[4649]=-76;
cos[4650]=-76;
cos[4651]=-76;
cos[4652]=-76;
cos[4653]=-76;
cos[4654]=-76;
cos[4655]=-76;
cos[4656]=-76;
cos[4657]=-76;
cos[4658]=-76;
cos[4659]=-76;
cos[4660]=-76;
cos[4661]=-76;
cos[4662]=-76;
cos[4663]=-76;
cos[4664]=-76;
cos[4665]=-76;
cos[4666]=-76;
cos[4667]=-76;
cos[4668]=-76;
cos[4669]=-76;
cos[4670]=-76;
cos[4671]=-76;
cos[4672]=-76;
cos[4673]=-76;
cos[4674]=-76;
cos[4675]=-77;
cos[4676]=-77;
cos[4677]=-77;
cos[4678]=-77;
cos[4679]=-77;
cos[4680]=-77;
cos[4681]=-77;
cos[4682]=-77;
cos[4683]=-77;
cos[4684]=-77;
cos[4685]=-77;
cos[4686]=-77;
cos[4687]=-77;
cos[4688]=-77;
cos[4689]=-77;
cos[4690]=-77;
cos[4691]=-77;
cos[4692]=-77;
cos[4693]=-77;
cos[4694]=-77;
cos[4695]=-77;
cos[4696]=-77;
cos[4697]=-77;
cos[4698]=-77;
cos[4699]=-77;
cos[4700]=-77;
cos[4701]=-77;
cos[4702]=-77;
cos[4703]=-77;
cos[4704]=-77;
cos[4705]=-77;
cos[4706]=-77;
cos[4707]=-77;
cos[4708]=-77;
cos[4709]=-77;
cos[4710]=-77;
cos[4711]=-77;
cos[4712]=-77;
cos[4713]=-77;
cos[4714]=-77;
cos[4715]=-77;
cos[4716]=-77;
cos[4717]=-77;
cos[4718]=-77;
cos[4719]=-77;
cos[4720]=-77;
cos[4721]=-77;
cos[4722]=-77;
cos[4723]=-77;
cos[4724]=-77;
cos[4725]=-77;
cos[4726]=-77;
cos[4727]=-77;
cos[4728]=-77;
cos[4729]=-77;
cos[4730]=-77;
cos[4731]=-77;
cos[4732]=-77;
cos[4733]=-77;
cos[4734]=-77;
cos[4735]=-77;
cos[4736]=-77;
cos[4737]=-77;
cos[4738]=-77;
cos[4739]=-77;
cos[4740]=-77;
cos[4741]=-77;
cos[4742]=-77;
cos[4743]=-77;
cos[4744]=-77;
cos[4745]=-77;
cos[4746]=-77;
cos[4747]=-77;
cos[4748]=-77;
cos[4749]=-77;
cos[4750]=-77;
cos[4751]=-77;
cos[4752]=-77;
cos[4753]=-77;
cos[4754]=-77;
cos[4755]=-77;
cos[4756]=-77;
cos[4757]=-77;
cos[4758]=-77;
cos[4759]=-77;
cos[4760]=-77;
cos[4761]=-77;
cos[4762]=-77;
cos[4763]=-77;
cos[4764]=-77;
cos[4765]=-77;
cos[4766]=-77;
cos[4767]=-77;
cos[4768]=-77;
cos[4769]=-77;
cos[4770]=-77;
cos[4771]=-77;
cos[4772]=-77;
cos[4773]=-77;
cos[4774]=-77;
cos[4775]=-77;
cos[4776]=-77;
cos[4777]=-77;
cos[4778]=-77;
cos[4779]=-77;
cos[4780]=-77;
cos[4781]=-77;
cos[4782]=-77;
cos[4783]=-77;
cos[4784]=-77;
cos[4785]=-77;
cos[4786]=-77;
cos[4787]=-77;
cos[4788]=-77;
cos[4789]=-77;
cos[4790]=-77;
cos[4791]=-77;
cos[4792]=-77;
cos[4793]=-77;
cos[4794]=-77;
cos[4795]=-77;
cos[4796]=-77;
cos[4797]=-77;
cos[4798]=-77;
cos[4799]=-78;
cos[4800]=-78;
cos[4801]=-78;
cos[4802]=-78;
cos[4803]=-78;
cos[4804]=-78;
cos[4805]=-78;
cos[4806]=-78;
cos[4807]=-78;
cos[4808]=-78;
cos[4809]=-78;
cos[4810]=-78;
cos[4811]=-78;
cos[4812]=-78;
cos[4813]=-78;
cos[4814]=-78;
cos[4815]=-78;
cos[4816]=-78;
cos[4817]=-78;
cos[4818]=-78;
cos[4819]=-78;
cos[4820]=-78;
cos[4821]=-78;
cos[4822]=-78;
cos[4823]=-78;
cos[4824]=-78;
cos[4825]=-78;
cos[4826]=-78;
cos[4827]=-78;
cos[4828]=-78;
cos[4829]=-78;
cos[4830]=-78;
cos[4831]=-78;
cos[4832]=-78;
cos[4833]=-78;
cos[4834]=-78;
cos[4835]=-78;
cos[4836]=-78;
cos[4837]=-78;
cos[4838]=-78;
cos[4839]=-78;
cos[4840]=-78;
cos[4841]=-78;
cos[4842]=-78;
cos[4843]=-78;
cos[4844]=-78;
cos[4845]=-78;
cos[4846]=-78;
cos[4847]=-78;
cos[4848]=-78;
cos[4849]=-78;
cos[4850]=-78;
cos[4851]=-78;
cos[4852]=-78;
cos[4853]=-78;
cos[4854]=-78;
cos[4855]=-78;
cos[4856]=-78;
cos[4857]=-78;
cos[4858]=-78;
cos[4859]=-78;
cos[4860]=-78;
cos[4861]=-78;
cos[4862]=-78;
cos[4863]=-78;
cos[4864]=-78;
cos[4865]=-78;
cos[4866]=-78;
cos[4867]=-78;
cos[4868]=-78;
cos[4869]=-78;
cos[4870]=-78;
cos[4871]=-78;
cos[4872]=-78;
cos[4873]=-78;
cos[4874]=-78;
cos[4875]=-78;
cos[4876]=-78;
cos[4877]=-78;
cos[4878]=-78;
cos[4879]=-78;
cos[4880]=-78;
cos[4881]=-78;
cos[4882]=-78;
cos[4883]=-78;
cos[4884]=-78;
cos[4885]=-78;
cos[4886]=-78;
cos[4887]=-78;
cos[4888]=-78;
cos[4889]=-78;
cos[4890]=-78;
cos[4891]=-78;
cos[4892]=-78;
cos[4893]=-78;
cos[4894]=-78;
cos[4895]=-78;
cos[4896]=-78;
cos[4897]=-78;
cos[4898]=-78;
cos[4899]=-78;
cos[4900]=-78;
cos[4901]=-78;
cos[4902]=-78;
cos[4903]=-78;
cos[4904]=-78;
cos[4905]=-78;
cos[4906]=-78;
cos[4907]=-78;
cos[4908]=-78;
cos[4909]=-78;
cos[4910]=-78;
cos[4911]=-78;
cos[4912]=-78;
cos[4913]=-78;
cos[4914]=-78;
cos[4915]=-78;
cos[4916]=-78;
cos[4917]=-78;
cos[4918]=-78;
cos[4919]=-78;
cos[4920]=-78;
cos[4921]=-78;
cos[4922]=-78;
cos[4923]=-78;
cos[4924]=-78;
cos[4925]=-78;
cos[4926]=-78;
cos[4927]=-78;
cos[4928]=-78;
cos[4929]=-78;
cos[4930]=-78;
cos[4931]=-78;
cos[4932]=-78;
cos[4933]=-78;
cos[4934]=-78;
cos[4935]=-78;
cos[4936]=-78;
cos[4937]=-78;
cos[4938]=-78;
cos[4939]=-78;
cos[4940]=-78;
cos[4941]=-78;
cos[4942]=-78;
cos[4943]=-78;
cos[4944]=-78;
cos[4945]=-78;
cos[4946]=-78;
cos[4947]=-78;
cos[4948]=-78;
cos[4949]=-78;
cos[4950]=-78;
cos[4951]=-78;
cos[4952]=-78;
cos[4953]=-78;
cos[4954]=-78;
cos[4955]=-78;
cos[4956]=-78;
cos[4957]=-78;
cos[4958]=-78;
cos[4959]=-78;
cos[4960]=-78;
cos[4961]=-78;
cos[4962]=-78;
cos[4963]=-78;
cos[4964]=-78;
cos[4965]=-78;
cos[4966]=-78;
cos[4967]=-78;
cos[4968]=-78;
cos[4969]=-78;
cos[4970]=-78;
cos[4971]=-78;
cos[4972]=-78;
cos[4973]=-78;
cos[4974]=-78;
cos[4975]=-78;
cos[4976]=-78;
cos[4977]=-78;
cos[4978]=-78;
cos[4979]=-78;
cos[4980]=-78;
cos[4981]=-78;
cos[4982]=-78;
cos[4983]=-78;
cos[4984]=-78;
cos[4985]=-78;
cos[4986]=-78;
cos[4987]=-78;
cos[4988]=-78;
cos[4989]=-78;
cos[4990]=-78;
cos[4991]=-78;
cos[4992]=-78;
cos[4993]=-78;
cos[4994]=-78;
cos[4995]=-78;
cos[4996]=-78;
cos[4997]=-78;
cos[4998]=-78;
cos[4999]=-78;
cos[5000]=-78;
cos[5001]=-78;
cos[5002]=-78;
cos[5003]=-78;
cos[5004]=-78;
cos[5005]=-78;
cos[5006]=-78;
cos[5007]=-78;
cos[5008]=-78;
cos[5009]=-78;
cos[5010]=-78;
cos[5011]=-78;
cos[5012]=-78;
cos[5013]=-78;
cos[5014]=-78;
cos[5015]=-78;
cos[5016]=-78;
cos[5017]=-78;
cos[5018]=-78;
cos[5019]=-78;
cos[5020]=-78;
cos[5021]=-78;
cos[5022]=-78;
cos[5023]=-78;
cos[5024]=-78;
cos[5025]=-78;
cos[5026]=-78;
cos[5027]=-78;
cos[5028]=-78;
cos[5029]=-78;
cos[5030]=-78;
cos[5031]=-78;
cos[5032]=-78;
cos[5033]=-78;
cos[5034]=-78;
cos[5035]=-78;
cos[5036]=-78;
cos[5037]=-78;
cos[5038]=-78;
cos[5039]=-78;
cos[5040]=-78;
cos[5041]=-78;
cos[5042]=-78;
cos[5043]=-78;
cos[5044]=-78;
cos[5045]=-78;
cos[5046]=-78;
cos[5047]=-78;
cos[5048]=-78;
cos[5049]=-78;
cos[5050]=-78;
cos[5051]=-78;
cos[5052]=-78;
cos[5053]=-78;
cos[5054]=-78;
cos[5055]=-78;
cos[5056]=-78;
cos[5057]=-78;
cos[5058]=-78;
cos[5059]=-78;
cos[5060]=-78;
cos[5061]=-78;
cos[5062]=-78;
cos[5063]=-78;
cos[5064]=-78;
cos[5065]=-78;
cos[5066]=-78;
cos[5067]=-78;
cos[5068]=-78;
cos[5069]=-78;
cos[5070]=-78;
cos[5071]=-78;
cos[5072]=-78;
cos[5073]=-78;
cos[5074]=-78;
cos[5075]=-78;
cos[5076]=-78;
cos[5077]=-78;
cos[5078]=-78;
cos[5079]=-78;
cos[5080]=-78;
cos[5081]=-78;
cos[5082]=-78;
cos[5083]=-78;
cos[5084]=-78;
cos[5085]=-78;
cos[5086]=-78;
cos[5087]=-78;
cos[5088]=-78;
cos[5089]=-78;
cos[5090]=-78;
cos[5091]=-78;
cos[5092]=-78;
cos[5093]=-78;
cos[5094]=-78;
cos[5095]=-78;
cos[5096]=-78;
cos[5097]=-78;
cos[5098]=-78;
cos[5099]=-78;
cos[5100]=-78;
cos[5101]=-78;
cos[5102]=-78;
cos[5103]=-78;
cos[5104]=-78;
cos[5105]=-78;
cos[5106]=-78;
cos[5107]=-78;
cos[5108]=-78;
cos[5109]=-78;
cos[5110]=-78;
cos[5111]=-78;
cos[5112]=-78;
cos[5113]=-78;
cos[5114]=-78;
cos[5115]=-78;
cos[5116]=-78;
cos[5117]=-78;
cos[5118]=-78;
cos[5119]=-78;
cos[5120]=-78;
cos[5121]=-78;
cos[5122]=-78;
cos[5123]=-78;
cos[5124]=-78;
cos[5125]=-78;
cos[5126]=-78;
cos[5127]=-78;
cos[5128]=-78;
cos[5129]=-78;
cos[5130]=-78;
cos[5131]=-78;
cos[5132]=-78;
cos[5133]=-78;
cos[5134]=-78;
cos[5135]=-78;
cos[5136]=-78;
cos[5137]=-78;
cos[5138]=-78;
cos[5139]=-78;
cos[5140]=-78;
cos[5141]=-78;
cos[5142]=-78;
cos[5143]=-78;
cos[5144]=-78;
cos[5145]=-78;
cos[5146]=-78;
cos[5147]=-78;
cos[5148]=-78;
cos[5149]=-78;
cos[5150]=-78;
cos[5151]=-78;
cos[5152]=-78;
cos[5153]=-78;
cos[5154]=-78;
cos[5155]=-78;
cos[5156]=-78;
cos[5157]=-78;
cos[5158]=-78;
cos[5159]=-78;
cos[5160]=-78;
cos[5161]=-78;
cos[5162]=-78;
cos[5163]=-78;
cos[5164]=-78;
cos[5165]=-78;
cos[5166]=-78;
cos[5167]=-78;
cos[5168]=-78;
cos[5169]=-78;
cos[5170]=-78;
cos[5171]=-78;
cos[5172]=-78;
cos[5173]=-78;
cos[5174]=-78;
cos[5175]=-78;
cos[5176]=-78;
cos[5177]=-78;
cos[5178]=-78;
cos[5179]=-78;
cos[5180]=-78;
cos[5181]=-78;
cos[5182]=-78;
cos[5183]=-78;
cos[5184]=-78;
cos[5185]=-78;
cos[5186]=-78;
cos[5187]=-78;
cos[5188]=-78;
cos[5189]=-78;
cos[5190]=-78;
cos[5191]=-78;
cos[5192]=-78;
cos[5193]=-78;
cos[5194]=-78;
cos[5195]=-78;
cos[5196]=-78;
cos[5197]=-78;
cos[5198]=-78;
cos[5199]=-78;
cos[5200]=-78;
cos[5201]=-78;
cos[5202]=-77;
cos[5203]=-77;
cos[5204]=-77;
cos[5205]=-77;
cos[5206]=-77;
cos[5207]=-77;
cos[5208]=-77;
cos[5209]=-77;
cos[5210]=-77;
cos[5211]=-77;
cos[5212]=-77;
cos[5213]=-77;
cos[5214]=-77;
cos[5215]=-77;
cos[5216]=-77;
cos[5217]=-77;
cos[5218]=-77;
cos[5219]=-77;
cos[5220]=-77;
cos[5221]=-77;
cos[5222]=-77;
cos[5223]=-77;
cos[5224]=-77;
cos[5225]=-77;
cos[5226]=-77;
cos[5227]=-77;
cos[5228]=-77;
cos[5229]=-77;
cos[5230]=-77;
cos[5231]=-77;
cos[5232]=-77;
cos[5233]=-77;
cos[5234]=-77;
cos[5235]=-77;
cos[5236]=-77;
cos[5237]=-77;
cos[5238]=-77;
cos[5239]=-77;
cos[5240]=-77;
cos[5241]=-77;
cos[5242]=-77;
cos[5243]=-77;
cos[5244]=-77;
cos[5245]=-77;
cos[5246]=-77;
cos[5247]=-77;
cos[5248]=-77;
cos[5249]=-77;
cos[5250]=-77;
cos[5251]=-77;
cos[5252]=-77;
cos[5253]=-77;
cos[5254]=-77;
cos[5255]=-77;
cos[5256]=-77;
cos[5257]=-77;
cos[5258]=-77;
cos[5259]=-77;
cos[5260]=-77;
cos[5261]=-77;
cos[5262]=-77;
cos[5263]=-77;
cos[5264]=-77;
cos[5265]=-77;
cos[5266]=-77;
cos[5267]=-77;
cos[5268]=-77;
cos[5269]=-77;
cos[5270]=-77;
cos[5271]=-77;
cos[5272]=-77;
cos[5273]=-77;
cos[5274]=-77;
cos[5275]=-77;
cos[5276]=-77;
cos[5277]=-77;
cos[5278]=-77;
cos[5279]=-77;
cos[5280]=-77;
cos[5281]=-77;
cos[5282]=-77;
cos[5283]=-77;
cos[5284]=-77;
cos[5285]=-77;
cos[5286]=-77;
cos[5287]=-77;
cos[5288]=-77;
cos[5289]=-77;
cos[5290]=-77;
cos[5291]=-77;
cos[5292]=-77;
cos[5293]=-77;
cos[5294]=-77;
cos[5295]=-77;
cos[5296]=-77;
cos[5297]=-77;
cos[5298]=-77;
cos[5299]=-77;
cos[5300]=-77;
cos[5301]=-77;
cos[5302]=-77;
cos[5303]=-77;
cos[5304]=-77;
cos[5305]=-77;
cos[5306]=-77;
cos[5307]=-77;
cos[5308]=-77;
cos[5309]=-77;
cos[5310]=-77;
cos[5311]=-77;
cos[5312]=-77;
cos[5313]=-77;
cos[5314]=-77;
cos[5315]=-77;
cos[5316]=-77;
cos[5317]=-77;
cos[5318]=-77;
cos[5319]=-77;
cos[5320]=-77;
cos[5321]=-77;
cos[5322]=-77;
cos[5323]=-77;
cos[5324]=-77;
cos[5325]=-77;
cos[5326]=-76;
cos[5327]=-76;
cos[5328]=-76;
cos[5329]=-76;
cos[5330]=-76;
cos[5331]=-76;
cos[5332]=-76;
cos[5333]=-76;
cos[5334]=-76;
cos[5335]=-76;
cos[5336]=-76;
cos[5337]=-76;
cos[5338]=-76;
cos[5339]=-76;
cos[5340]=-76;
cos[5341]=-76;
cos[5342]=-76;
cos[5343]=-76;
cos[5344]=-76;
cos[5345]=-76;
cos[5346]=-76;
cos[5347]=-76;
cos[5348]=-76;
cos[5349]=-76;
cos[5350]=-76;
cos[5351]=-76;
cos[5352]=-76;
cos[5353]=-76;
cos[5354]=-76;
cos[5355]=-76;
cos[5356]=-76;
cos[5357]=-76;
cos[5358]=-76;
cos[5359]=-76;
cos[5360]=-76;
cos[5361]=-76;
cos[5362]=-76;
cos[5363]=-76;
cos[5364]=-76;
cos[5365]=-76;
cos[5366]=-76;
cos[5367]=-76;
cos[5368]=-76;
cos[5369]=-76;
cos[5370]=-76;
cos[5371]=-76;
cos[5372]=-76;
cos[5373]=-76;
cos[5374]=-76;
cos[5375]=-76;
cos[5376]=-76;
cos[5377]=-76;
cos[5378]=-76;
cos[5379]=-76;
cos[5380]=-76;
cos[5381]=-76;
cos[5382]=-76;
cos[5383]=-76;
cos[5384]=-76;
cos[5385]=-76;
cos[5386]=-76;
cos[5387]=-76;
cos[5388]=-76;
cos[5389]=-76;
cos[5390]=-76;
cos[5391]=-76;
cos[5392]=-76;
cos[5393]=-76;
cos[5394]=-76;
cos[5395]=-76;
cos[5396]=-76;
cos[5397]=-76;
cos[5398]=-76;
cos[5399]=-76;
cos[5400]=-76;
cos[5401]=-76;
cos[5402]=-76;
cos[5403]=-76;
cos[5404]=-76;
cos[5405]=-76;
cos[5406]=-76;
cos[5407]=-76;
cos[5408]=-76;
cos[5409]=-76;
cos[5410]=-76;
cos[5411]=-76;
cos[5412]=-76;
cos[5413]=-76;
cos[5414]=-75;
cos[5415]=-75;
cos[5416]=-75;
cos[5417]=-75;
cos[5418]=-75;
cos[5419]=-75;
cos[5420]=-75;
cos[5421]=-75;
cos[5422]=-75;
cos[5423]=-75;
cos[5424]=-75;
cos[5425]=-75;
cos[5426]=-75;
cos[5427]=-75;
cos[5428]=-75;
cos[5429]=-75;
cos[5430]=-75;
cos[5431]=-75;
cos[5432]=-75;
cos[5433]=-75;
cos[5434]=-75;
cos[5435]=-75;
cos[5436]=-75;
cos[5437]=-75;
cos[5438]=-75;
cos[5439]=-75;
cos[5440]=-75;
cos[5441]=-75;
cos[5442]=-75;
cos[5443]=-75;
cos[5444]=-75;
cos[5445]=-75;
cos[5446]=-75;
cos[5447]=-75;
cos[5448]=-75;
cos[5449]=-75;
cos[5450]=-75;
cos[5451]=-75;
cos[5452]=-75;
cos[5453]=-75;
cos[5454]=-75;
cos[5455]=-75;
cos[5456]=-75;
cos[5457]=-75;
cos[5458]=-75;
cos[5459]=-75;
cos[5460]=-75;
cos[5461]=-75;
cos[5462]=-75;
cos[5463]=-75;
cos[5464]=-75;
cos[5465]=-75;
cos[5466]=-75;
cos[5467]=-75;
cos[5468]=-75;
cos[5469]=-75;
cos[5470]=-75;
cos[5471]=-75;
cos[5472]=-75;
cos[5473]=-75;
cos[5474]=-75;
cos[5475]=-75;
cos[5476]=-75;
cos[5477]=-75;
cos[5478]=-75;
cos[5479]=-75;
cos[5480]=-75;
cos[5481]=-75;
cos[5482]=-75;
cos[5483]=-75;
cos[5484]=-75;
cos[5485]=-75;
cos[5486]=-75;
cos[5487]=-74;
cos[5488]=-74;
cos[5489]=-74;
cos[5490]=-74;
cos[5491]=-74;
cos[5492]=-74;
cos[5493]=-74;
cos[5494]=-74;
cos[5495]=-74;
cos[5496]=-74;
cos[5497]=-74;
cos[5498]=-74;
cos[5499]=-74;
cos[5500]=-74;
cos[5501]=-74;
cos[5502]=-74;
cos[5503]=-74;
cos[5504]=-74;
cos[5505]=-74;
cos[5506]=-74;
cos[5507]=-74;
cos[5508]=-74;
cos[5509]=-74;
cos[5510]=-74;
cos[5511]=-74;
cos[5512]=-74;
cos[5513]=-74;
cos[5514]=-74;
cos[5515]=-74;
cos[5516]=-74;
cos[5517]=-74;
cos[5518]=-74;
cos[5519]=-74;
cos[5520]=-74;
cos[5521]=-74;
cos[5522]=-74;
cos[5523]=-74;
cos[5524]=-74;
cos[5525]=-74;
cos[5526]=-74;
cos[5527]=-74;
cos[5528]=-74;
cos[5529]=-74;
cos[5530]=-74;
cos[5531]=-74;
cos[5532]=-74;
cos[5533]=-74;
cos[5534]=-74;
cos[5535]=-74;
cos[5536]=-74;
cos[5537]=-74;
cos[5538]=-74;
cos[5539]=-74;
cos[5540]=-74;
cos[5541]=-74;
cos[5542]=-74;
cos[5543]=-74;
cos[5544]=-74;
cos[5545]=-74;
cos[5546]=-74;
cos[5547]=-74;
cos[5548]=-74;
cos[5549]=-74;
cos[5550]=-74;
cos[5551]=-73;
cos[5552]=-73;
cos[5553]=-73;
cos[5554]=-73;
cos[5555]=-73;
cos[5556]=-73;
cos[5557]=-73;
cos[5558]=-73;
cos[5559]=-73;
cos[5560]=-73;
cos[5561]=-73;
cos[5562]=-73;
cos[5563]=-73;
cos[5564]=-73;
cos[5565]=-73;
cos[5566]=-73;
cos[5567]=-73;
cos[5568]=-73;
cos[5569]=-73;
cos[5570]=-73;
cos[5571]=-73;
cos[5572]=-73;
cos[5573]=-73;
cos[5574]=-73;
cos[5575]=-73;
cos[5576]=-73;
cos[5577]=-73;
cos[5578]=-73;
cos[5579]=-73;
cos[5580]=-73;
cos[5581]=-73;
cos[5582]=-73;
cos[5583]=-73;
cos[5584]=-73;
cos[5585]=-73;
cos[5586]=-73;
cos[5587]=-73;
cos[5588]=-73;
cos[5589]=-73;
cos[5590]=-73;
cos[5591]=-73;
cos[5592]=-73;
cos[5593]=-73;
cos[5594]=-73;
cos[5595]=-73;
cos[5596]=-73;
cos[5597]=-73;
cos[5598]=-73;
cos[5599]=-73;
cos[5600]=-73;
cos[5601]=-73;
cos[5602]=-73;
cos[5603]=-73;
cos[5604]=-73;
cos[5605]=-73;
cos[5606]=-73;
cos[5607]=-73;
cos[5608]=-72;
cos[5609]=-72;
cos[5610]=-72;
cos[5611]=-72;
cos[5612]=-72;
cos[5613]=-72;
cos[5614]=-72;
cos[5615]=-72;
cos[5616]=-72;
cos[5617]=-72;
cos[5618]=-72;
cos[5619]=-72;
cos[5620]=-72;
cos[5621]=-72;
cos[5622]=-72;
cos[5623]=-72;
cos[5624]=-72;
cos[5625]=-72;
cos[5626]=-72;
cos[5627]=-72;
cos[5628]=-72;
cos[5629]=-72;
cos[5630]=-72;
cos[5631]=-72;
cos[5632]=-72;
cos[5633]=-72;
cos[5634]=-72;
cos[5635]=-72;
cos[5636]=-72;
cos[5637]=-72;
cos[5638]=-72;
cos[5639]=-72;
cos[5640]=-72;
cos[5641]=-72;
cos[5642]=-72;
cos[5643]=-72;
cos[5644]=-72;
cos[5645]=-72;
cos[5646]=-72;
cos[5647]=-72;
cos[5648]=-72;
cos[5649]=-72;
cos[5650]=-72;
cos[5651]=-72;
cos[5652]=-72;
cos[5653]=-72;
cos[5654]=-72;
cos[5655]=-72;
cos[5656]=-72;
cos[5657]=-72;
cos[5658]=-72;
cos[5659]=-72;
cos[5660]=-72;
cos[5661]=-71;
cos[5662]=-71;
cos[5663]=-71;
cos[5664]=-71;
cos[5665]=-71;
cos[5666]=-71;
cos[5667]=-71;
cos[5668]=-71;
cos[5669]=-71;
cos[5670]=-71;
cos[5671]=-71;
cos[5672]=-71;
cos[5673]=-71;
cos[5674]=-71;
cos[5675]=-71;
cos[5676]=-71;
cos[5677]=-71;
cos[5678]=-71;
cos[5679]=-71;
cos[5680]=-71;
cos[5681]=-71;
cos[5682]=-71;
cos[5683]=-71;
cos[5684]=-71;
cos[5685]=-71;
cos[5686]=-71;
cos[5687]=-71;
cos[5688]=-71;
cos[5689]=-71;
cos[5690]=-71;
cos[5691]=-71;
cos[5692]=-71;
cos[5693]=-71;
cos[5694]=-71;
cos[5695]=-71;
cos[5696]=-71;
cos[5697]=-71;
cos[5698]=-71;
cos[5699]=-71;
cos[5700]=-71;
cos[5701]=-71;
cos[5702]=-71;
cos[5703]=-71;
cos[5704]=-71;
cos[5705]=-71;
cos[5706]=-71;
cos[5707]=-71;
cos[5708]=-71;
cos[5709]=-71;
cos[5710]=-70;
cos[5711]=-70;
cos[5712]=-70;
cos[5713]=-70;
cos[5714]=-70;
cos[5715]=-70;
cos[5716]=-70;
cos[5717]=-70;
cos[5718]=-70;
cos[5719]=-70;
cos[5720]=-70;
cos[5721]=-70;
cos[5722]=-70;
cos[5723]=-70;
cos[5724]=-70;
cos[5725]=-70;
cos[5726]=-70;
cos[5727]=-70;
cos[5728]=-70;
cos[5729]=-70;
cos[5730]=-70;
cos[5731]=-70;
cos[5732]=-70;
cos[5733]=-70;
cos[5734]=-70;
cos[5735]=-70;
cos[5736]=-70;
cos[5737]=-70;
cos[5738]=-70;
cos[5739]=-70;
cos[5740]=-70;
cos[5741]=-70;
cos[5742]=-70;
cos[5743]=-70;
cos[5744]=-70;
cos[5745]=-70;
cos[5746]=-70;
cos[5747]=-70;
cos[5748]=-70;
cos[5749]=-70;
cos[5750]=-70;
cos[5751]=-70;
cos[5752]=-70;
cos[5753]=-70;
cos[5754]=-70;
cos[5755]=-69;
cos[5756]=-69;
cos[5757]=-69;
cos[5758]=-69;
cos[5759]=-69;
cos[5760]=-69;
cos[5761]=-69;
cos[5762]=-69;
cos[5763]=-69;
cos[5764]=-69;
cos[5765]=-69;
cos[5766]=-69;
cos[5767]=-69;
cos[5768]=-69;
cos[5769]=-69;
cos[5770]=-69;
cos[5771]=-69;
cos[5772]=-69;
cos[5773]=-69;
cos[5774]=-69;
cos[5775]=-69;
cos[5776]=-69;
cos[5777]=-69;
cos[5778]=-69;
cos[5779]=-69;
cos[5780]=-69;
cos[5781]=-69;
cos[5782]=-69;
cos[5783]=-69;
cos[5784]=-69;
cos[5785]=-69;
cos[5786]=-69;
cos[5787]=-69;
cos[5788]=-69;
cos[5789]=-69;
cos[5790]=-69;
cos[5791]=-69;
cos[5792]=-69;
cos[5793]=-69;
cos[5794]=-69;
cos[5795]=-69;
cos[5796]=-69;
cos[5797]=-69;
cos[5798]=-69;
cos[5799]=-68;
cos[5800]=-68;
cos[5801]=-68;
cos[5802]=-68;
cos[5803]=-68;
cos[5804]=-68;
cos[5805]=-68;
cos[5806]=-68;
cos[5807]=-68;
cos[5808]=-68;
cos[5809]=-68;
cos[5810]=-68;
cos[5811]=-68;
cos[5812]=-68;
cos[5813]=-68;
cos[5814]=-68;
cos[5815]=-68;
cos[5816]=-68;
cos[5817]=-68;
cos[5818]=-68;
cos[5819]=-68;
cos[5820]=-68;
cos[5821]=-68;
cos[5822]=-68;
cos[5823]=-68;
cos[5824]=-68;
cos[5825]=-68;
cos[5826]=-68;
cos[5827]=-68;
cos[5828]=-68;
cos[5829]=-68;
cos[5830]=-68;
cos[5831]=-68;
cos[5832]=-68;
cos[5833]=-68;
cos[5834]=-68;
cos[5835]=-68;
cos[5836]=-68;
cos[5837]=-68;
cos[5838]=-68;
cos[5839]=-68;
cos[5840]=-67;
cos[5841]=-67;
cos[5842]=-67;
cos[5843]=-67;
cos[5844]=-67;
cos[5845]=-67;
cos[5846]=-67;
cos[5847]=-67;
cos[5848]=-67;
cos[5849]=-67;
cos[5850]=-67;
cos[5851]=-67;
cos[5852]=-67;
cos[5853]=-67;
cos[5854]=-67;
cos[5855]=-67;
cos[5856]=-67;
cos[5857]=-67;
cos[5858]=-67;
cos[5859]=-67;
cos[5860]=-67;
cos[5861]=-67;
cos[5862]=-67;
cos[5863]=-67;
cos[5864]=-67;
cos[5865]=-67;
cos[5866]=-67;
cos[5867]=-67;
cos[5868]=-67;
cos[5869]=-67;
cos[5870]=-67;
cos[5871]=-67;
cos[5872]=-67;
cos[5873]=-67;
cos[5874]=-67;
cos[5875]=-67;
cos[5876]=-67;
cos[5877]=-67;
cos[5878]=-67;
cos[5879]=-67;
cos[5880]=-66;
cos[5881]=-66;
cos[5882]=-66;
cos[5883]=-66;
cos[5884]=-66;
cos[5885]=-66;
cos[5886]=-66;
cos[5887]=-66;
cos[5888]=-66;
cos[5889]=-66;
cos[5890]=-66;
cos[5891]=-66;
cos[5892]=-66;
cos[5893]=-66;
cos[5894]=-66;
cos[5895]=-66;
cos[5896]=-66;
cos[5897]=-66;
cos[5898]=-66;
cos[5899]=-66;
cos[5900]=-66;
cos[5901]=-66;
cos[5902]=-66;
cos[5903]=-66;
cos[5904]=-66;
cos[5905]=-66;
cos[5906]=-66;
cos[5907]=-66;
cos[5908]=-66;
cos[5909]=-66;
cos[5910]=-66;
cos[5911]=-66;
cos[5912]=-66;
cos[5913]=-66;
cos[5914]=-66;
cos[5915]=-66;
cos[5916]=-66;
cos[5917]=-66;
cos[5918]=-65;
cos[5919]=-65;
cos[5920]=-65;
cos[5921]=-65;
cos[5922]=-65;
cos[5923]=-65;
cos[5924]=-65;
cos[5925]=-65;
cos[5926]=-65;
cos[5927]=-65;
cos[5928]=-65;
cos[5929]=-65;
cos[5930]=-65;
cos[5931]=-65;
cos[5932]=-65;
cos[5933]=-65;
cos[5934]=-65;
cos[5935]=-65;
cos[5936]=-65;
cos[5937]=-65;
cos[5938]=-65;
cos[5939]=-65;
cos[5940]=-65;
cos[5941]=-65;
cos[5942]=-65;
cos[5943]=-65;
cos[5944]=-65;
cos[5945]=-65;
cos[5946]=-65;
cos[5947]=-65;
cos[5948]=-65;
cos[5949]=-65;
cos[5950]=-65;
cos[5951]=-65;
cos[5952]=-65;
cos[5953]=-65;
cos[5954]=-65;
cos[5955]=-64;
cos[5956]=-64;
cos[5957]=-64;
cos[5958]=-64;
cos[5959]=-64;
cos[5960]=-64;
cos[5961]=-64;
cos[5962]=-64;
cos[5963]=-64;
cos[5964]=-64;
cos[5965]=-64;
cos[5966]=-64;
cos[5967]=-64;
cos[5968]=-64;
cos[5969]=-64;
cos[5970]=-64;
cos[5971]=-64;
cos[5972]=-64;
cos[5973]=-64;
cos[5974]=-64;
cos[5975]=-64;
cos[5976]=-64;
cos[5977]=-64;
cos[5978]=-64;
cos[5979]=-64;
cos[5980]=-64;
cos[5981]=-64;
cos[5982]=-64;
cos[5983]=-64;
cos[5984]=-64;
cos[5985]=-64;
cos[5986]=-64;
cos[5987]=-64;
cos[5988]=-64;
cos[5989]=-64;
cos[5990]=-63;
cos[5991]=-63;
cos[5992]=-63;
cos[5993]=-63;
cos[5994]=-63;
cos[5995]=-63;
cos[5996]=-63;
cos[5997]=-63;
cos[5998]=-63;
cos[5999]=-63;
cos[6000]=-63;
cos[6001]=-63;
cos[6002]=-63;
cos[6003]=-63;
cos[6004]=-63;
cos[6005]=-63;
cos[6006]=-63;
cos[6007]=-63;
cos[6008]=-63;
cos[6009]=-63;
cos[6010]=-63;
cos[6011]=-63;
cos[6012]=-63;
cos[6013]=-63;
cos[6014]=-63;
cos[6015]=-63;
cos[6016]=-63;
cos[6017]=-63;
cos[6018]=-63;
cos[6019]=-63;
cos[6020]=-63;
cos[6021]=-63;
cos[6022]=-63;
cos[6023]=-63;
cos[6024]=-63;
cos[6025]=-62;
cos[6026]=-62;
cos[6027]=-62;
cos[6028]=-62;
cos[6029]=-62;
cos[6030]=-62;
cos[6031]=-62;
cos[6032]=-62;
cos[6033]=-62;
cos[6034]=-62;
cos[6035]=-62;
cos[6036]=-62;
cos[6037]=-62;
cos[6038]=-62;
cos[6039]=-62;
cos[6040]=-62;
cos[6041]=-62;
cos[6042]=-62;
cos[6043]=-62;
cos[6044]=-62;
cos[6045]=-62;
cos[6046]=-62;
cos[6047]=-62;
cos[6048]=-62;
cos[6049]=-62;
cos[6050]=-62;
cos[6051]=-62;
cos[6052]=-62;
cos[6053]=-62;
cos[6054]=-62;
cos[6055]=-62;
cos[6056]=-62;
cos[6057]=-62;
cos[6058]=-61;
cos[6059]=-61;
cos[6060]=-61;
cos[6061]=-61;
cos[6062]=-61;
cos[6063]=-61;
cos[6064]=-61;
cos[6065]=-61;
cos[6066]=-61;
cos[6067]=-61;
cos[6068]=-61;
cos[6069]=-61;
cos[6070]=-61;
cos[6071]=-61;
cos[6072]=-61;
cos[6073]=-61;
cos[6074]=-61;
cos[6075]=-61;
cos[6076]=-61;
cos[6077]=-61;
cos[6078]=-61;
cos[6079]=-61;
cos[6080]=-61;
cos[6081]=-61;
cos[6082]=-61;
cos[6083]=-61;
cos[6084]=-61;
cos[6085]=-61;
cos[6086]=-61;
cos[6087]=-61;
cos[6088]=-61;
cos[6089]=-61;
cos[6090]=-61;
cos[6091]=-60;
cos[6092]=-60;
cos[6093]=-60;
cos[6094]=-60;
cos[6095]=-60;
cos[6096]=-60;
cos[6097]=-60;
cos[6098]=-60;
cos[6099]=-60;
cos[6100]=-60;
cos[6101]=-60;
cos[6102]=-60;
cos[6103]=-60;
cos[6104]=-60;
cos[6105]=-60;
cos[6106]=-60;
cos[6107]=-60;
cos[6108]=-60;
cos[6109]=-60;
cos[6110]=-60;
cos[6111]=-60;
cos[6112]=-60;
cos[6113]=-60;
cos[6114]=-60;
cos[6115]=-60;
cos[6116]=-60;
cos[6117]=-60;
cos[6118]=-60;
cos[6119]=-60;
cos[6120]=-60;
cos[6121]=-60;
cos[6122]=-60;
cos[6123]=-59;
cos[6124]=-59;
cos[6125]=-59;
cos[6126]=-59;
cos[6127]=-59;
cos[6128]=-59;
cos[6129]=-59;
cos[6130]=-59;
cos[6131]=-59;
cos[6132]=-59;
cos[6133]=-59;
cos[6134]=-59;
cos[6135]=-59;
cos[6136]=-59;
cos[6137]=-59;
cos[6138]=-59;
cos[6139]=-59;
cos[6140]=-59;
cos[6141]=-59;
cos[6142]=-59;
cos[6143]=-59;
cos[6144]=-59;
cos[6145]=-59;
cos[6146]=-59;
cos[6147]=-59;
cos[6148]=-59;
cos[6149]=-59;
cos[6150]=-59;
cos[6151]=-59;
cos[6152]=-59;
cos[6153]=-59;
cos[6154]=-58;
cos[6155]=-58;
cos[6156]=-58;
cos[6157]=-58;
cos[6158]=-58;
cos[6159]=-58;
cos[6160]=-58;
cos[6161]=-58;
cos[6162]=-58;
cos[6163]=-58;
cos[6164]=-58;
cos[6165]=-58;
cos[6166]=-58;
cos[6167]=-58;
cos[6168]=-58;
cos[6169]=-58;
cos[6170]=-58;
cos[6171]=-58;
cos[6172]=-58;
cos[6173]=-58;
cos[6174]=-58;
cos[6175]=-58;
cos[6176]=-58;
cos[6177]=-58;
cos[6178]=-58;
cos[6179]=-58;
cos[6180]=-58;
cos[6181]=-58;
cos[6182]=-58;
cos[6183]=-58;
cos[6184]=-57;
cos[6185]=-57;
cos[6186]=-57;
cos[6187]=-57;
cos[6188]=-57;
cos[6189]=-57;
cos[6190]=-57;
cos[6191]=-57;
cos[6192]=-57;
cos[6193]=-57;
cos[6194]=-57;
cos[6195]=-57;
cos[6196]=-57;
cos[6197]=-57;
cos[6198]=-57;
cos[6199]=-57;
cos[6200]=-57;
cos[6201]=-57;
cos[6202]=-57;
cos[6203]=-57;
cos[6204]=-57;
cos[6205]=-57;
cos[6206]=-57;
cos[6207]=-57;
cos[6208]=-57;
cos[6209]=-57;
cos[6210]=-57;
cos[6211]=-57;
cos[6212]=-57;
cos[6213]=-57;
cos[6214]=-56;
cos[6215]=-56;
cos[6216]=-56;
cos[6217]=-56;
cos[6218]=-56;
cos[6219]=-56;
cos[6220]=-56;
cos[6221]=-56;
cos[6222]=-56;
cos[6223]=-56;
cos[6224]=-56;
cos[6225]=-56;
cos[6226]=-56;
cos[6227]=-56;
cos[6228]=-56;
cos[6229]=-56;
cos[6230]=-56;
cos[6231]=-56;
cos[6232]=-56;
cos[6233]=-56;
cos[6234]=-56;
cos[6235]=-56;
cos[6236]=-56;
cos[6237]=-56;
cos[6238]=-56;
cos[6239]=-56;
cos[6240]=-56;
cos[6241]=-56;
cos[6242]=-56;
cos[6243]=-55;
cos[6244]=-55;
cos[6245]=-55;
cos[6246]=-55;
cos[6247]=-55;
cos[6248]=-55;
cos[6249]=-55;
cos[6250]=-55;
cos[6251]=-55;
cos[6252]=-55;
cos[6253]=-55;
cos[6254]=-55;
cos[6255]=-55;
cos[6256]=-55;
cos[6257]=-55;
cos[6258]=-55;
cos[6259]=-55;
cos[6260]=-55;
cos[6261]=-55;
cos[6262]=-55;
cos[6263]=-55;
cos[6264]=-55;
cos[6265]=-55;
cos[6266]=-55;
cos[6267]=-55;
cos[6268]=-55;
cos[6269]=-55;
cos[6270]=-55;
cos[6271]=-55;
cos[6272]=-54;
cos[6273]=-54;
cos[6274]=-54;
cos[6275]=-54;
cos[6276]=-54;
cos[6277]=-54;
cos[6278]=-54;
cos[6279]=-54;
cos[6280]=-54;
cos[6281]=-54;
cos[6282]=-54;
cos[6283]=-54;
cos[6284]=-54;
cos[6285]=-54;
cos[6286]=-54;
cos[6287]=-54;
cos[6288]=-54;
cos[6289]=-54;
cos[6290]=-54;
cos[6291]=-54;
cos[6292]=-54;
cos[6293]=-54;
cos[6294]=-54;
cos[6295]=-54;
cos[6296]=-54;
cos[6297]=-54;
cos[6298]=-54;
cos[6299]=-54;
cos[6300]=-53;
cos[6301]=-53;
cos[6302]=-53;
cos[6303]=-53;
cos[6304]=-53;
cos[6305]=-53;
cos[6306]=-53;
cos[6307]=-53;
cos[6308]=-53;
cos[6309]=-53;
cos[6310]=-53;
cos[6311]=-53;
cos[6312]=-53;
cos[6313]=-53;
cos[6314]=-53;
cos[6315]=-53;
cos[6316]=-53;
cos[6317]=-53;
cos[6318]=-53;
cos[6319]=-53;
cos[6320]=-53;
cos[6321]=-53;
cos[6322]=-53;
cos[6323]=-53;
cos[6324]=-53;
cos[6325]=-53;
cos[6326]=-53;
cos[6327]=-53;
cos[6328]=-52;
cos[6329]=-52;
cos[6330]=-52;
cos[6331]=-52;
cos[6332]=-52;
cos[6333]=-52;
cos[6334]=-52;
cos[6335]=-52;
cos[6336]=-52;
cos[6337]=-52;
cos[6338]=-52;
cos[6339]=-52;
cos[6340]=-52;
cos[6341]=-52;
cos[6342]=-52;
cos[6343]=-52;
cos[6344]=-52;
cos[6345]=-52;
cos[6346]=-52;
cos[6347]=-52;
cos[6348]=-52;
cos[6349]=-52;
cos[6350]=-52;
cos[6351]=-52;
cos[6352]=-52;
cos[6353]=-52;
cos[6354]=-52;
cos[6355]=-51;
cos[6356]=-51;
cos[6357]=-51;
cos[6358]=-51;
cos[6359]=-51;
cos[6360]=-51;
cos[6361]=-51;
cos[6362]=-51;
cos[6363]=-51;
cos[6364]=-51;
cos[6365]=-51;
cos[6366]=-51;
cos[6367]=-51;
cos[6368]=-51;
cos[6369]=-51;
cos[6370]=-51;
cos[6371]=-51;
cos[6372]=-51;
cos[6373]=-51;
cos[6374]=-51;
cos[6375]=-51;
cos[6376]=-51;
cos[6377]=-51;
cos[6378]=-51;
cos[6379]=-51;
cos[6380]=-51;
cos[6381]=-51;
cos[6382]=-50;
cos[6383]=-50;
cos[6384]=-50;
cos[6385]=-50;
cos[6386]=-50;
cos[6387]=-50;
cos[6388]=-50;
cos[6389]=-50;
cos[6390]=-50;
cos[6391]=-50;
cos[6392]=-50;
cos[6393]=-50;
cos[6394]=-50;
cos[6395]=-50;
cos[6396]=-50;
cos[6397]=-50;
cos[6398]=-50;
cos[6399]=-50;
cos[6400]=-50;
cos[6401]=-50;
cos[6402]=-50;
cos[6403]=-50;
cos[6404]=-50;
cos[6405]=-50;
cos[6406]=-50;
cos[6407]=-50;
cos[6408]=-49;
cos[6409]=-49;
cos[6410]=-49;
cos[6411]=-49;
cos[6412]=-49;
cos[6413]=-49;
cos[6414]=-49;
cos[6415]=-49;
cos[6416]=-49;
cos[6417]=-49;
cos[6418]=-49;
cos[6419]=-49;
cos[6420]=-49;
cos[6421]=-49;
cos[6422]=-49;
cos[6423]=-49;
cos[6424]=-49;
cos[6425]=-49;
cos[6426]=-49;
cos[6427]=-49;
cos[6428]=-49;
cos[6429]=-49;
cos[6430]=-49;
cos[6431]=-49;
cos[6432]=-49;
cos[6433]=-49;
cos[6434]=-49;
cos[6435]=-48;
cos[6436]=-48;
cos[6437]=-48;
cos[6438]=-48;
cos[6439]=-48;
cos[6440]=-48;
cos[6441]=-48;
cos[6442]=-48;
cos[6443]=-48;
cos[6444]=-48;
cos[6445]=-48;
cos[6446]=-48;
cos[6447]=-48;
cos[6448]=-48;
cos[6449]=-48;
cos[6450]=-48;
cos[6451]=-48;
cos[6452]=-48;
cos[6453]=-48;
cos[6454]=-48;
cos[6455]=-48;
cos[6456]=-48;
cos[6457]=-48;
cos[6458]=-48;
cos[6459]=-48;
cos[6460]=-47;
cos[6461]=-47;
cos[6462]=-47;
cos[6463]=-47;
cos[6464]=-47;
cos[6465]=-47;
cos[6466]=-47;
cos[6467]=-47;
cos[6468]=-47;
cos[6469]=-47;
cos[6470]=-47;
cos[6471]=-47;
cos[6472]=-47;
cos[6473]=-47;
cos[6474]=-47;
cos[6475]=-47;
cos[6476]=-47;
cos[6477]=-47;
cos[6478]=-47;
cos[6479]=-47;
cos[6480]=-47;
cos[6481]=-47;
cos[6482]=-47;
cos[6483]=-47;
cos[6484]=-47;
cos[6485]=-47;
cos[6486]=-46;
cos[6487]=-46;
cos[6488]=-46;
cos[6489]=-46;
cos[6490]=-46;
cos[6491]=-46;
cos[6492]=-46;
cos[6493]=-46;
cos[6494]=-46;
cos[6495]=-46;
cos[6496]=-46;
cos[6497]=-46;
cos[6498]=-46;
cos[6499]=-46;
cos[6500]=-46;
cos[6501]=-46;
cos[6502]=-46;
cos[6503]=-46;
cos[6504]=-46;
cos[6505]=-46;
cos[6506]=-46;
cos[6507]=-46;
cos[6508]=-46;
cos[6509]=-46;
cos[6510]=-46;
cos[6511]=-45;
cos[6512]=-45;
cos[6513]=-45;
cos[6514]=-45;
cos[6515]=-45;
cos[6516]=-45;
cos[6517]=-45;
cos[6518]=-45;
cos[6519]=-45;
cos[6520]=-45;
cos[6521]=-45;
cos[6522]=-45;
cos[6523]=-45;
cos[6524]=-45;
cos[6525]=-45;
cos[6526]=-45;
cos[6527]=-45;
cos[6528]=-45;
cos[6529]=-45;
cos[6530]=-45;
cos[6531]=-45;
cos[6532]=-45;
cos[6533]=-45;
cos[6534]=-45;
cos[6535]=-45;
cos[6536]=-44;
cos[6537]=-44;
cos[6538]=-44;
cos[6539]=-44;
cos[6540]=-44;
cos[6541]=-44;
cos[6542]=-44;
cos[6543]=-44;
cos[6544]=-44;
cos[6545]=-44;
cos[6546]=-44;
cos[6547]=-44;
cos[6548]=-44;
cos[6549]=-44;
cos[6550]=-44;
cos[6551]=-44;
cos[6552]=-44;
cos[6553]=-44;
cos[6554]=-44;
cos[6555]=-44;
cos[6556]=-44;
cos[6557]=-44;
cos[6558]=-44;
cos[6559]=-44;
cos[6560]=-44;
cos[6561]=-43;
cos[6562]=-43;
cos[6563]=-43;
cos[6564]=-43;
cos[6565]=-43;
cos[6566]=-43;
cos[6567]=-43;
cos[6568]=-43;
cos[6569]=-43;
cos[6570]=-43;
cos[6571]=-43;
cos[6572]=-43;
cos[6573]=-43;
cos[6574]=-43;
cos[6575]=-43;
cos[6576]=-43;
cos[6577]=-43;
cos[6578]=-43;
cos[6579]=-43;
cos[6580]=-43;
cos[6581]=-43;
cos[6582]=-43;
cos[6583]=-43;
cos[6584]=-43;
cos[6585]=-42;
cos[6586]=-42;
cos[6587]=-42;
cos[6588]=-42;
cos[6589]=-42;
cos[6590]=-42;
cos[6591]=-42;
cos[6592]=-42;
cos[6593]=-42;
cos[6594]=-42;
cos[6595]=-42;
cos[6596]=-42;
cos[6597]=-42;
cos[6598]=-42;
cos[6599]=-42;
cos[6600]=-42;
cos[6601]=-42;
cos[6602]=-42;
cos[6603]=-42;
cos[6604]=-42;
cos[6605]=-42;
cos[6606]=-42;
cos[6607]=-42;
cos[6608]=-42;
cos[6609]=-41;
cos[6610]=-41;
cos[6611]=-41;
cos[6612]=-41;
cos[6613]=-41;
cos[6614]=-41;
cos[6615]=-41;
cos[6616]=-41;
cos[6617]=-41;
cos[6618]=-41;
cos[6619]=-41;
cos[6620]=-41;
cos[6621]=-41;
cos[6622]=-41;
cos[6623]=-41;
cos[6624]=-41;
cos[6625]=-41;
cos[6626]=-41;
cos[6627]=-41;
cos[6628]=-41;
cos[6629]=-41;
cos[6630]=-41;
cos[6631]=-41;
cos[6632]=-41;
cos[6633]=-40;
cos[6634]=-40;
cos[6635]=-40;
cos[6636]=-40;
cos[6637]=-40;
cos[6638]=-40;
cos[6639]=-40;
cos[6640]=-40;
cos[6641]=-40;
cos[6642]=-40;
cos[6643]=-40;
cos[6644]=-40;
cos[6645]=-40;
cos[6646]=-40;
cos[6647]=-40;
cos[6648]=-40;
cos[6649]=-40;
cos[6650]=-40;
cos[6651]=-40;
cos[6652]=-40;
cos[6653]=-40;
cos[6654]=-40;
cos[6655]=-40;
cos[6656]=-40;
cos[6657]=-39;
cos[6658]=-39;
cos[6659]=-39;
cos[6660]=-39;
cos[6661]=-39;
cos[6662]=-39;
cos[6663]=-39;
cos[6664]=-39;
cos[6665]=-39;
cos[6666]=-39;
cos[6667]=-39;
cos[6668]=-39;
cos[6669]=-39;
cos[6670]=-39;
cos[6671]=-39;
cos[6672]=-39;
cos[6673]=-39;
cos[6674]=-39;
cos[6675]=-39;
cos[6676]=-39;
cos[6677]=-39;
cos[6678]=-39;
cos[6679]=-39;
cos[6680]=-38;
cos[6681]=-38;
cos[6682]=-38;
cos[6683]=-38;
cos[6684]=-38;
cos[6685]=-38;
cos[6686]=-38;
cos[6687]=-38;
cos[6688]=-38;
cos[6689]=-38;
cos[6690]=-38;
cos[6691]=-38;
cos[6692]=-38;
cos[6693]=-38;
cos[6694]=-38;
cos[6695]=-38;
cos[6696]=-38;
cos[6697]=-38;
cos[6698]=-38;
cos[6699]=-38;
cos[6700]=-38;
cos[6701]=-38;
cos[6702]=-38;
cos[6703]=-38;
cos[6704]=-37;
cos[6705]=-37;
cos[6706]=-37;
cos[6707]=-37;
cos[6708]=-37;
cos[6709]=-37;
cos[6710]=-37;
cos[6711]=-37;
cos[6712]=-37;
cos[6713]=-37;
cos[6714]=-37;
cos[6715]=-37;
cos[6716]=-37;
cos[6717]=-37;
cos[6718]=-37;
cos[6719]=-37;
cos[6720]=-37;
cos[6721]=-37;
cos[6722]=-37;
cos[6723]=-37;
cos[6724]=-37;
cos[6725]=-37;
cos[6726]=-37;
cos[6727]=-36;
cos[6728]=-36;
cos[6729]=-36;
cos[6730]=-36;
cos[6731]=-36;
cos[6732]=-36;
cos[6733]=-36;
cos[6734]=-36;
cos[6735]=-36;
cos[6736]=-36;
cos[6737]=-36;
cos[6738]=-36;
cos[6739]=-36;
cos[6740]=-36;
cos[6741]=-36;
cos[6742]=-36;
cos[6743]=-36;
cos[6744]=-36;
cos[6745]=-36;
cos[6746]=-36;
cos[6747]=-36;
cos[6748]=-36;
cos[6749]=-36;
cos[6750]=-35;
cos[6751]=-35;
cos[6752]=-35;
cos[6753]=-35;
cos[6754]=-35;
cos[6755]=-35;
cos[6756]=-35;
cos[6757]=-35;
cos[6758]=-35;
cos[6759]=-35;
cos[6760]=-35;
cos[6761]=-35;
cos[6762]=-35;
cos[6763]=-35;
cos[6764]=-35;
cos[6765]=-35;
cos[6766]=-35;
cos[6767]=-35;
cos[6768]=-35;
cos[6769]=-35;
cos[6770]=-35;
cos[6771]=-35;
cos[6772]=-35;
cos[6773]=-34;
cos[6774]=-34;
cos[6775]=-34;
cos[6776]=-34;
cos[6777]=-34;
cos[6778]=-34;
cos[6779]=-34;
cos[6780]=-34;
cos[6781]=-34;
cos[6782]=-34;
cos[6783]=-34;
cos[6784]=-34;
cos[6785]=-34;
cos[6786]=-34;
cos[6787]=-34;
cos[6788]=-34;
cos[6789]=-34;
cos[6790]=-34;
cos[6791]=-34;
cos[6792]=-34;
cos[6793]=-34;
cos[6794]=-34;
cos[6795]=-33;
cos[6796]=-33;
cos[6797]=-33;
cos[6798]=-33;
cos[6799]=-33;
cos[6800]=-33;
cos[6801]=-33;
cos[6802]=-33;
cos[6803]=-33;
cos[6804]=-33;
cos[6805]=-33;
cos[6806]=-33;
cos[6807]=-33;
cos[6808]=-33;
cos[6809]=-33;
cos[6810]=-33;
cos[6811]=-33;
cos[6812]=-33;
cos[6813]=-33;
cos[6814]=-33;
cos[6815]=-33;
cos[6816]=-33;
cos[6817]=-33;
cos[6818]=-32;
cos[6819]=-32;
cos[6820]=-32;
cos[6821]=-32;
cos[6822]=-32;
cos[6823]=-32;
cos[6824]=-32;
cos[6825]=-32;
cos[6826]=-32;
cos[6827]=-32;
cos[6828]=-32;
cos[6829]=-32;
cos[6830]=-32;
cos[6831]=-32;
cos[6832]=-32;
cos[6833]=-32;
cos[6834]=-32;
cos[6835]=-32;
cos[6836]=-32;
cos[6837]=-32;
cos[6838]=-32;
cos[6839]=-32;
cos[6840]=-31;
cos[6841]=-31;
cos[6842]=-31;
cos[6843]=-31;
cos[6844]=-31;
cos[6845]=-31;
cos[6846]=-31;
cos[6847]=-31;
cos[6848]=-31;
cos[6849]=-31;
cos[6850]=-31;
cos[6851]=-31;
cos[6852]=-31;
cos[6853]=-31;
cos[6854]=-31;
cos[6855]=-31;
cos[6856]=-31;
cos[6857]=-31;
cos[6858]=-31;
cos[6859]=-31;
cos[6860]=-31;
cos[6861]=-31;
cos[6862]=-30;
cos[6863]=-30;
cos[6864]=-30;
cos[6865]=-30;
cos[6866]=-30;
cos[6867]=-30;
cos[6868]=-30;
cos[6869]=-30;
cos[6870]=-30;
cos[6871]=-30;
cos[6872]=-30;
cos[6873]=-30;
cos[6874]=-30;
cos[6875]=-30;
cos[6876]=-30;
cos[6877]=-30;
cos[6878]=-30;
cos[6879]=-30;
cos[6880]=-30;
cos[6881]=-30;
cos[6882]=-30;
cos[6883]=-30;
cos[6884]=-29;
cos[6885]=-29;
cos[6886]=-29;
cos[6887]=-29;
cos[6888]=-29;
cos[6889]=-29;
cos[6890]=-29;
cos[6891]=-29;
cos[6892]=-29;
cos[6893]=-29;
cos[6894]=-29;
cos[6895]=-29;
cos[6896]=-29;
cos[6897]=-29;
cos[6898]=-29;
cos[6899]=-29;
cos[6900]=-29;
cos[6901]=-29;
cos[6902]=-29;
cos[6903]=-29;
cos[6904]=-29;
cos[6905]=-29;
cos[6906]=-28;
cos[6907]=-28;
cos[6908]=-28;
cos[6909]=-28;
cos[6910]=-28;
cos[6911]=-28;
cos[6912]=-28;
cos[6913]=-28;
cos[6914]=-28;
cos[6915]=-28;
cos[6916]=-28;
cos[6917]=-28;
cos[6918]=-28;
cos[6919]=-28;
cos[6920]=-28;
cos[6921]=-28;
cos[6922]=-28;
cos[6923]=-28;
cos[6924]=-28;
cos[6925]=-28;
cos[6926]=-28;
cos[6927]=-28;
cos[6928]=-27;
cos[6929]=-27;
cos[6930]=-27;
cos[6931]=-27;
cos[6932]=-27;
cos[6933]=-27;
cos[6934]=-27;
cos[6935]=-27;
cos[6936]=-27;
cos[6937]=-27;
cos[6938]=-27;
cos[6939]=-27;
cos[6940]=-27;
cos[6941]=-27;
cos[6942]=-27;
cos[6943]=-27;
cos[6944]=-27;
cos[6945]=-27;
cos[6946]=-27;
cos[6947]=-27;
cos[6948]=-27;
cos[6949]=-27;
cos[6950]=-26;
cos[6951]=-26;
cos[6952]=-26;
cos[6953]=-26;
cos[6954]=-26;
cos[6955]=-26;
cos[6956]=-26;
cos[6957]=-26;
cos[6958]=-26;
cos[6959]=-26;
cos[6960]=-26;
cos[6961]=-26;
cos[6962]=-26;
cos[6963]=-26;
cos[6964]=-26;
cos[6965]=-26;
cos[6966]=-26;
cos[6967]=-26;
cos[6968]=-26;
cos[6969]=-26;
cos[6970]=-26;
cos[6971]=-25;
cos[6972]=-25;
cos[6973]=-25;
cos[6974]=-25;
cos[6975]=-25;
cos[6976]=-25;
cos[6977]=-25;
cos[6978]=-25;
cos[6979]=-25;
cos[6980]=-25;
cos[6981]=-25;
cos[6982]=-25;
cos[6983]=-25;
cos[6984]=-25;
cos[6985]=-25;
cos[6986]=-25;
cos[6987]=-25;
cos[6988]=-25;
cos[6989]=-25;
cos[6990]=-25;
cos[6991]=-25;
cos[6992]=-25;
cos[6993]=-24;
cos[6994]=-24;
cos[6995]=-24;
cos[6996]=-24;
cos[6997]=-24;
cos[6998]=-24;
cos[6999]=-24;
cos[7000]=-24;
cos[7001]=-24;
cos[7002]=-24;
cos[7003]=-24;
cos[7004]=-24;
cos[7005]=-24;
cos[7006]=-24;
cos[7007]=-24;
cos[7008]=-24;
cos[7009]=-24;
cos[7010]=-24;
cos[7011]=-24;
cos[7012]=-24;
cos[7013]=-24;
cos[7014]=-23;
cos[7015]=-23;
cos[7016]=-23;
cos[7017]=-23;
cos[7018]=-23;
cos[7019]=-23;
cos[7020]=-23;
cos[7021]=-23;
cos[7022]=-23;
cos[7023]=-23;
cos[7024]=-23;
cos[7025]=-23;
cos[7026]=-23;
cos[7027]=-23;
cos[7028]=-23;
cos[7029]=-23;
cos[7030]=-23;
cos[7031]=-23;
cos[7032]=-23;
cos[7033]=-23;
cos[7034]=-23;
cos[7035]=-23;
cos[7036]=-22;
cos[7037]=-22;
cos[7038]=-22;
cos[7039]=-22;
cos[7040]=-22;
cos[7041]=-22;
cos[7042]=-22;
cos[7043]=-22;
cos[7044]=-22;
cos[7045]=-22;
cos[7046]=-22;
cos[7047]=-22;
cos[7048]=-22;
cos[7049]=-22;
cos[7050]=-22;
cos[7051]=-22;
cos[7052]=-22;
cos[7053]=-22;
cos[7054]=-22;
cos[7055]=-22;
cos[7056]=-22;
cos[7057]=-21;
cos[7058]=-21;
cos[7059]=-21;
cos[7060]=-21;
cos[7061]=-21;
cos[7062]=-21;
cos[7063]=-21;
cos[7064]=-21;
cos[7065]=-21;
cos[7066]=-21;
cos[7067]=-21;
cos[7068]=-21;
cos[7069]=-21;
cos[7070]=-21;
cos[7071]=-21;
cos[7072]=-21;
cos[7073]=-21;
cos[7074]=-21;
cos[7075]=-21;
cos[7076]=-21;
cos[7077]=-21;
cos[7078]=-20;
cos[7079]=-20;
cos[7080]=-20;
cos[7081]=-20;
cos[7082]=-20;
cos[7083]=-20;
cos[7084]=-20;
cos[7085]=-20;
cos[7086]=-20;
cos[7087]=-20;
cos[7088]=-20;
cos[7089]=-20;
cos[7090]=-20;
cos[7091]=-20;
cos[7092]=-20;
cos[7093]=-20;
cos[7094]=-20;
cos[7095]=-20;
cos[7096]=-20;
cos[7097]=-20;
cos[7098]=-20;
cos[7099]=-19;
cos[7100]=-19;
cos[7101]=-19;
cos[7102]=-19;
cos[7103]=-19;
cos[7104]=-19;
cos[7105]=-19;
cos[7106]=-19;
cos[7107]=-19;
cos[7108]=-19;
cos[7109]=-19;
cos[7110]=-19;
cos[7111]=-19;
cos[7112]=-19;
cos[7113]=-19;
cos[7114]=-19;
cos[7115]=-19;
cos[7116]=-19;
cos[7117]=-19;
cos[7118]=-19;
cos[7119]=-19;
cos[7120]=-18;
cos[7121]=-18;
cos[7122]=-18;
cos[7123]=-18;
cos[7124]=-18;
cos[7125]=-18;
cos[7126]=-18;
cos[7127]=-18;
cos[7128]=-18;
cos[7129]=-18;
cos[7130]=-18;
cos[7131]=-18;
cos[7132]=-18;
cos[7133]=-18;
cos[7134]=-18;
cos[7135]=-18;
cos[7136]=-18;
cos[7137]=-18;
cos[7138]=-18;
cos[7139]=-18;
cos[7140]=-18;
cos[7141]=-17;
cos[7142]=-17;
cos[7143]=-17;
cos[7144]=-17;
cos[7145]=-17;
cos[7146]=-17;
cos[7147]=-17;
cos[7148]=-17;
cos[7149]=-17;
cos[7150]=-17;
cos[7151]=-17;
cos[7152]=-17;
cos[7153]=-17;
cos[7154]=-17;
cos[7155]=-17;
cos[7156]=-17;
cos[7157]=-17;
cos[7158]=-17;
cos[7159]=-17;
cos[7160]=-17;
cos[7161]=-17;
cos[7162]=-16;
cos[7163]=-16;
cos[7164]=-16;
cos[7165]=-16;
cos[7166]=-16;
cos[7167]=-16;
cos[7168]=-16;
cos[7169]=-16;
cos[7170]=-16;
cos[7171]=-16;
cos[7172]=-16;
cos[7173]=-16;
cos[7174]=-16;
cos[7175]=-16;
cos[7176]=-16;
cos[7177]=-16;
cos[7178]=-16;
cos[7179]=-16;
cos[7180]=-16;
cos[7181]=-16;
cos[7182]=-16;
cos[7183]=-15;
cos[7184]=-15;
cos[7185]=-15;
cos[7186]=-15;
cos[7187]=-15;
cos[7188]=-15;
cos[7189]=-15;
cos[7190]=-15;
cos[7191]=-15;
cos[7192]=-15;
cos[7193]=-15;
cos[7194]=-15;
cos[7195]=-15;
cos[7196]=-15;
cos[7197]=-15;
cos[7198]=-15;
cos[7199]=-15;
cos[7200]=-15;
cos[7201]=-15;
cos[7202]=-15;
cos[7203]=-14;
cos[7204]=-14;
cos[7205]=-14;
cos[7206]=-14;
cos[7207]=-14;
cos[7208]=-14;
cos[7209]=-14;
cos[7210]=-14;
cos[7211]=-14;
cos[7212]=-14;
cos[7213]=-14;
cos[7214]=-14;
cos[7215]=-14;
cos[7216]=-14;
cos[7217]=-14;
cos[7218]=-14;
cos[7219]=-14;
cos[7220]=-14;
cos[7221]=-14;
cos[7222]=-14;
cos[7223]=-14;
cos[7224]=-13;
cos[7225]=-13;
cos[7226]=-13;
cos[7227]=-13;
cos[7228]=-13;
cos[7229]=-13;
cos[7230]=-13;
cos[7231]=-13;
cos[7232]=-13;
cos[7233]=-13;
cos[7234]=-13;
cos[7235]=-13;
cos[7236]=-13;
cos[7237]=-13;
cos[7238]=-13;
cos[7239]=-13;
cos[7240]=-13;
cos[7241]=-13;
cos[7242]=-13;
cos[7243]=-13;
cos[7244]=-13;
cos[7245]=-12;
cos[7246]=-12;
cos[7247]=-12;
cos[7248]=-12;
cos[7249]=-12;
cos[7250]=-12;
cos[7251]=-12;
cos[7252]=-12;
cos[7253]=-12;
cos[7254]=-12;
cos[7255]=-12;
cos[7256]=-12;
cos[7257]=-12;
cos[7258]=-12;
cos[7259]=-12;
cos[7260]=-12;
cos[7261]=-12;
cos[7262]=-12;
cos[7263]=-12;
cos[7264]=-12;
cos[7265]=-11;
cos[7266]=-11;
cos[7267]=-11;
cos[7268]=-11;
cos[7269]=-11;
cos[7270]=-11;
cos[7271]=-11;
cos[7272]=-11;
cos[7273]=-11;
cos[7274]=-11;
cos[7275]=-11;
cos[7276]=-11;
cos[7277]=-11;
cos[7278]=-11;
cos[7279]=-11;
cos[7280]=-11;
cos[7281]=-11;
cos[7282]=-11;
cos[7283]=-11;
cos[7284]=-11;
cos[7285]=-11;
cos[7286]=-10;
cos[7287]=-10;
cos[7288]=-10;
cos[7289]=-10;
cos[7290]=-10;
cos[7291]=-10;
cos[7292]=-10;
cos[7293]=-10;
cos[7294]=-10;
cos[7295]=-10;
cos[7296]=-10;
cos[7297]=-10;
cos[7298]=-10;
cos[7299]=-10;
cos[7300]=-10;
cos[7301]=-10;
cos[7302]=-10;
cos[7303]=-10;
cos[7304]=-10;
cos[7305]=-10;
cos[7306]=-9;
cos[7307]=-9;
cos[7308]=-9;
cos[7309]=-9;
cos[7310]=-9;
cos[7311]=-9;
cos[7312]=-9;
cos[7313]=-9;
cos[7314]=-9;
cos[7315]=-9;
cos[7316]=-9;
cos[7317]=-9;
cos[7318]=-9;
cos[7319]=-9;
cos[7320]=-9;
cos[7321]=-9;
cos[7322]=-9;
cos[7323]=-9;
cos[7324]=-9;
cos[7325]=-9;
cos[7326]=-9;
cos[7327]=-8;
cos[7328]=-8;
cos[7329]=-8;
cos[7330]=-8;
cos[7331]=-8;
cos[7332]=-8;
cos[7333]=-8;
cos[7334]=-8;
cos[7335]=-8;
cos[7336]=-8;
cos[7337]=-8;
cos[7338]=-8;
cos[7339]=-8;
cos[7340]=-8;
cos[7341]=-8;
cos[7342]=-8;
cos[7343]=-8;
cos[7344]=-8;
cos[7345]=-8;
cos[7346]=-8;
cos[7347]=-7;
cos[7348]=-7;
cos[7349]=-7;
cos[7350]=-7;
cos[7351]=-7;
cos[7352]=-7;
cos[7353]=-7;
cos[7354]=-7;
cos[7355]=-7;
cos[7356]=-7;
cos[7357]=-7;
cos[7358]=-7;
cos[7359]=-7;
cos[7360]=-7;
cos[7361]=-7;
cos[7362]=-7;
cos[7363]=-7;
cos[7364]=-7;
cos[7365]=-7;
cos[7366]=-7;
cos[7367]=-7;
cos[7368]=-6;
cos[7369]=-6;
cos[7370]=-6;
cos[7371]=-6;
cos[7372]=-6;
cos[7373]=-6;
cos[7374]=-6;
cos[7375]=-6;
cos[7376]=-6;
cos[7377]=-6;
cos[7378]=-6;
cos[7379]=-6;
cos[7380]=-6;
cos[7381]=-6;
cos[7382]=-6;
cos[7383]=-6;
cos[7384]=-6;
cos[7385]=-6;
cos[7386]=-6;
cos[7387]=-6;
cos[7388]=-5;
cos[7389]=-5;
cos[7390]=-5;
cos[7391]=-5;
cos[7392]=-5;
cos[7393]=-5;
cos[7394]=-5;
cos[7395]=-5;
cos[7396]=-5;
cos[7397]=-5;
cos[7398]=-5;
cos[7399]=-5;
cos[7400]=-5;
cos[7401]=-5;
cos[7402]=-5;
cos[7403]=-5;
cos[7404]=-5;
cos[7405]=-5;
cos[7406]=-5;
cos[7407]=-5;
cos[7408]=-5;
cos[7409]=-4;
cos[7410]=-4;
cos[7411]=-4;
cos[7412]=-4;
cos[7413]=-4;
cos[7414]=-4;
cos[7415]=-4;
cos[7416]=-4;
cos[7417]=-4;
cos[7418]=-4;
cos[7419]=-4;
cos[7420]=-4;
cos[7421]=-4;
cos[7422]=-4;
cos[7423]=-4;
cos[7424]=-4;
cos[7425]=-4;
cos[7426]=-4;
cos[7427]=-4;
cos[7428]=-4;
cos[7429]=-3;
cos[7430]=-3;
cos[7431]=-3;
cos[7432]=-3;
cos[7433]=-3;
cos[7434]=-3;
cos[7435]=-3;
cos[7436]=-3;
cos[7437]=-3;
cos[7438]=-3;
cos[7439]=-3;
cos[7440]=-3;
cos[7441]=-3;
cos[7442]=-3;
cos[7443]=-3;
cos[7444]=-3;
cos[7445]=-3;
cos[7446]=-3;
cos[7447]=-3;
cos[7448]=-3;
cos[7449]=-3;
cos[7450]=-2;
cos[7451]=-2;
cos[7452]=-2;
cos[7453]=-2;
cos[7454]=-2;
cos[7455]=-2;
cos[7456]=-2;
cos[7457]=-2;
cos[7458]=-2;
cos[7459]=-2;
cos[7460]=-2;
cos[7461]=-2;
cos[7462]=-2;
cos[7463]=-2;
cos[7464]=-2;
cos[7465]=-2;
cos[7466]=-2;
cos[7467]=-2;
cos[7468]=-2;
cos[7469]=-2;
cos[7470]=-1;
cos[7471]=-1;
cos[7472]=-1;
cos[7473]=-1;
cos[7474]=-1;
cos[7475]=-1;
cos[7476]=-1;
cos[7477]=-1;
cos[7478]=-1;
cos[7479]=-1;
cos[7480]=-1;
cos[7481]=-1;
cos[7482]=-1;
cos[7483]=-1;
cos[7484]=-1;
cos[7485]=-1;
cos[7486]=-1;
cos[7487]=-1;
cos[7488]=-1;
cos[7489]=-1;
cos[7490]=0;
cos[7491]=0;
cos[7492]=0;
cos[7493]=0;
cos[7494]=0;
cos[7495]=0;
cos[7496]=0;
cos[7497]=0;
cos[7498]=0;
cos[7499]=0;
cos[7500]=0;
cos[7501]=0;
cos[7502]=0;
cos[7503]=0;
cos[7504]=0;
cos[7505]=0;
cos[7506]=0;
cos[7507]=0;
cos[7508]=0;
cos[7509]=0;
cos[7510]=0;
cos[7511]=1;
cos[7512]=1;
cos[7513]=1;
cos[7514]=1;
cos[7515]=1;
cos[7516]=1;
cos[7517]=1;
cos[7518]=1;
cos[7519]=1;
cos[7520]=1;
cos[7521]=1;
cos[7522]=1;
cos[7523]=1;
cos[7524]=1;
cos[7525]=1;
cos[7526]=1;
cos[7527]=1;
cos[7528]=1;
cos[7529]=1;
cos[7530]=1;
cos[7531]=2;
cos[7532]=2;
cos[7533]=2;
cos[7534]=2;
cos[7535]=2;
cos[7536]=2;
cos[7537]=2;
cos[7538]=2;
cos[7539]=2;
cos[7540]=2;
cos[7541]=2;
cos[7542]=2;
cos[7543]=2;
cos[7544]=2;
cos[7545]=2;
cos[7546]=2;
cos[7547]=2;
cos[7548]=2;
cos[7549]=2;
cos[7550]=2;
cos[7551]=3;
cos[7552]=3;
cos[7553]=3;
cos[7554]=3;
cos[7555]=3;
cos[7556]=3;
cos[7557]=3;
cos[7558]=3;
cos[7559]=3;
cos[7560]=3;
cos[7561]=3;
cos[7562]=3;
cos[7563]=3;
cos[7564]=3;
cos[7565]=3;
cos[7566]=3;
cos[7567]=3;
cos[7568]=3;
cos[7569]=3;
cos[7570]=3;
cos[7571]=3;
cos[7572]=4;
cos[7573]=4;
cos[7574]=4;
cos[7575]=4;
cos[7576]=4;
cos[7577]=4;
cos[7578]=4;
cos[7579]=4;
cos[7580]=4;
cos[7581]=4;
cos[7582]=4;
cos[7583]=4;
cos[7584]=4;
cos[7585]=4;
cos[7586]=4;
cos[7587]=4;
cos[7588]=4;
cos[7589]=4;
cos[7590]=4;
cos[7591]=4;
cos[7592]=5;
cos[7593]=5;
cos[7594]=5;
cos[7595]=5;
cos[7596]=5;
cos[7597]=5;
cos[7598]=5;
cos[7599]=5;
cos[7600]=5;
cos[7601]=5;
cos[7602]=5;
cos[7603]=5;
cos[7604]=5;
cos[7605]=5;
cos[7606]=5;
cos[7607]=5;
cos[7608]=5;
cos[7609]=5;
cos[7610]=5;
cos[7611]=5;
cos[7612]=5;
cos[7613]=6;
cos[7614]=6;
cos[7615]=6;
cos[7616]=6;
cos[7617]=6;
cos[7618]=6;
cos[7619]=6;
cos[7620]=6;
cos[7621]=6;
cos[7622]=6;
cos[7623]=6;
cos[7624]=6;
cos[7625]=6;
cos[7626]=6;
cos[7627]=6;
cos[7628]=6;
cos[7629]=6;
cos[7630]=6;
cos[7631]=6;
cos[7632]=6;
cos[7633]=7;
cos[7634]=7;
cos[7635]=7;
cos[7636]=7;
cos[7637]=7;
cos[7638]=7;
cos[7639]=7;
cos[7640]=7;
cos[7641]=7;
cos[7642]=7;
cos[7643]=7;
cos[7644]=7;
cos[7645]=7;
cos[7646]=7;
cos[7647]=7;
cos[7648]=7;
cos[7649]=7;
cos[7650]=7;
cos[7651]=7;
cos[7652]=7;
cos[7653]=7;
cos[7654]=8;
cos[7655]=8;
cos[7656]=8;
cos[7657]=8;
cos[7658]=8;
cos[7659]=8;
cos[7660]=8;
cos[7661]=8;
cos[7662]=8;
cos[7663]=8;
cos[7664]=8;
cos[7665]=8;
cos[7666]=8;
cos[7667]=8;
cos[7668]=8;
cos[7669]=8;
cos[7670]=8;
cos[7671]=8;
cos[7672]=8;
cos[7673]=8;
cos[7674]=9;
cos[7675]=9;
cos[7676]=9;
cos[7677]=9;
cos[7678]=9;
cos[7679]=9;
cos[7680]=9;
cos[7681]=9;
cos[7682]=9;
cos[7683]=9;
cos[7684]=9;
cos[7685]=9;
cos[7686]=9;
cos[7687]=9;
cos[7688]=9;
cos[7689]=9;
cos[7690]=9;
cos[7691]=9;
cos[7692]=9;
cos[7693]=9;
cos[7694]=9;
cos[7695]=10;
cos[7696]=10;
cos[7697]=10;
cos[7698]=10;
cos[7699]=10;
cos[7700]=10;
cos[7701]=10;
cos[7702]=10;
cos[7703]=10;
cos[7704]=10;
cos[7705]=10;
cos[7706]=10;
cos[7707]=10;
cos[7708]=10;
cos[7709]=10;
cos[7710]=10;
cos[7711]=10;
cos[7712]=10;
cos[7713]=10;
cos[7714]=10;
cos[7715]=11;
cos[7716]=11;
cos[7717]=11;
cos[7718]=11;
cos[7719]=11;
cos[7720]=11;
cos[7721]=11;
cos[7722]=11;
cos[7723]=11;
cos[7724]=11;
cos[7725]=11;
cos[7726]=11;
cos[7727]=11;
cos[7728]=11;
cos[7729]=11;
cos[7730]=11;
cos[7731]=11;
cos[7732]=11;
cos[7733]=11;
cos[7734]=11;
cos[7735]=11;
cos[7736]=12;
cos[7737]=12;
cos[7738]=12;
cos[7739]=12;
cos[7740]=12;
cos[7741]=12;
cos[7742]=12;
cos[7743]=12;
cos[7744]=12;
cos[7745]=12;
cos[7746]=12;
cos[7747]=12;
cos[7748]=12;
cos[7749]=12;
cos[7750]=12;
cos[7751]=12;
cos[7752]=12;
cos[7753]=12;
cos[7754]=12;
cos[7755]=12;
cos[7756]=13;
cos[7757]=13;
cos[7758]=13;
cos[7759]=13;
cos[7760]=13;
cos[7761]=13;
cos[7762]=13;
cos[7763]=13;
cos[7764]=13;
cos[7765]=13;
cos[7766]=13;
cos[7767]=13;
cos[7768]=13;
cos[7769]=13;
cos[7770]=13;
cos[7771]=13;
cos[7772]=13;
cos[7773]=13;
cos[7774]=13;
cos[7775]=13;
cos[7776]=13;
cos[7777]=14;
cos[7778]=14;
cos[7779]=14;
cos[7780]=14;
cos[7781]=14;
cos[7782]=14;
cos[7783]=14;
cos[7784]=14;
cos[7785]=14;
cos[7786]=14;
cos[7787]=14;
cos[7788]=14;
cos[7789]=14;
cos[7790]=14;
cos[7791]=14;
cos[7792]=14;
cos[7793]=14;
cos[7794]=14;
cos[7795]=14;
cos[7796]=14;
cos[7797]=14;
cos[7798]=15;
cos[7799]=15;
cos[7800]=15;
cos[7801]=15;
cos[7802]=15;
cos[7803]=15;
cos[7804]=15;
cos[7805]=15;
cos[7806]=15;
cos[7807]=15;
cos[7808]=15;
cos[7809]=15;
cos[7810]=15;
cos[7811]=15;
cos[7812]=15;
cos[7813]=15;
cos[7814]=15;
cos[7815]=15;
cos[7816]=15;
cos[7817]=15;
cos[7818]=16;
cos[7819]=16;
cos[7820]=16;
cos[7821]=16;
cos[7822]=16;
cos[7823]=16;
cos[7824]=16;
cos[7825]=16;
cos[7826]=16;
cos[7827]=16;
cos[7828]=16;
cos[7829]=16;
cos[7830]=16;
cos[7831]=16;
cos[7832]=16;
cos[7833]=16;
cos[7834]=16;
cos[7835]=16;
cos[7836]=16;
cos[7837]=16;
cos[7838]=16;
cos[7839]=17;
cos[7840]=17;
cos[7841]=17;
cos[7842]=17;
cos[7843]=17;
cos[7844]=17;
cos[7845]=17;
cos[7846]=17;
cos[7847]=17;
cos[7848]=17;
cos[7849]=17;
cos[7850]=17;
cos[7851]=17;
cos[7852]=17;
cos[7853]=17;
cos[7854]=17;
cos[7855]=17;
cos[7856]=17;
cos[7857]=17;
cos[7858]=17;
cos[7859]=17;
cos[7860]=18;
cos[7861]=18;
cos[7862]=18;
cos[7863]=18;
cos[7864]=18;
cos[7865]=18;
cos[7866]=18;
cos[7867]=18;
cos[7868]=18;
cos[7869]=18;
cos[7870]=18;
cos[7871]=18;
cos[7872]=18;
cos[7873]=18;
cos[7874]=18;
cos[7875]=18;
cos[7876]=18;
cos[7877]=18;
cos[7878]=18;
cos[7879]=18;
cos[7880]=18;
cos[7881]=19;
cos[7882]=19;
cos[7883]=19;
cos[7884]=19;
cos[7885]=19;
cos[7886]=19;
cos[7887]=19;
cos[7888]=19;
cos[7889]=19;
cos[7890]=19;
cos[7891]=19;
cos[7892]=19;
cos[7893]=19;
cos[7894]=19;
cos[7895]=19;
cos[7896]=19;
cos[7897]=19;
cos[7898]=19;
cos[7899]=19;
cos[7900]=19;
cos[7901]=19;
cos[7902]=20;
cos[7903]=20;
cos[7904]=20;
cos[7905]=20;
cos[7906]=20;
cos[7907]=20;
cos[7908]=20;
cos[7909]=20;
cos[7910]=20;
cos[7911]=20;
cos[7912]=20;
cos[7913]=20;
cos[7914]=20;
cos[7915]=20;
cos[7916]=20;
cos[7917]=20;
cos[7918]=20;
cos[7919]=20;
cos[7920]=20;
cos[7921]=20;
cos[7922]=20;
cos[7923]=21;
cos[7924]=21;
cos[7925]=21;
cos[7926]=21;
cos[7927]=21;
cos[7928]=21;
cos[7929]=21;
cos[7930]=21;
cos[7931]=21;
cos[7932]=21;
cos[7933]=21;
cos[7934]=21;
cos[7935]=21;
cos[7936]=21;
cos[7937]=21;
cos[7938]=21;
cos[7939]=21;
cos[7940]=21;
cos[7941]=21;
cos[7942]=21;
cos[7943]=21;
cos[7944]=22;
cos[7945]=22;
cos[7946]=22;
cos[7947]=22;
cos[7948]=22;
cos[7949]=22;
cos[7950]=22;
cos[7951]=22;
cos[7952]=22;
cos[7953]=22;
cos[7954]=22;
cos[7955]=22;
cos[7956]=22;
cos[7957]=22;
cos[7958]=22;
cos[7959]=22;
cos[7960]=22;
cos[7961]=22;
cos[7962]=22;
cos[7963]=22;
cos[7964]=22;
cos[7965]=23;
cos[7966]=23;
cos[7967]=23;
cos[7968]=23;
cos[7969]=23;
cos[7970]=23;
cos[7971]=23;
cos[7972]=23;
cos[7973]=23;
cos[7974]=23;
cos[7975]=23;
cos[7976]=23;
cos[7977]=23;
cos[7978]=23;
cos[7979]=23;
cos[7980]=23;
cos[7981]=23;
cos[7982]=23;
cos[7983]=23;
cos[7984]=23;
cos[7985]=23;
cos[7986]=23;
cos[7987]=24;
cos[7988]=24;
cos[7989]=24;
cos[7990]=24;
cos[7991]=24;
cos[7992]=24;
cos[7993]=24;
cos[7994]=24;
cos[7995]=24;
cos[7996]=24;
cos[7997]=24;
cos[7998]=24;
cos[7999]=24;
cos[8000]=24;
cos[8001]=24;
cos[8002]=24;
cos[8003]=24;
cos[8004]=24;
cos[8005]=24;
cos[8006]=24;
cos[8007]=24;
cos[8008]=25;
cos[8009]=25;
cos[8010]=25;
cos[8011]=25;
cos[8012]=25;
cos[8013]=25;
cos[8014]=25;
cos[8015]=25;
cos[8016]=25;
cos[8017]=25;
cos[8018]=25;
cos[8019]=25;
cos[8020]=25;
cos[8021]=25;
cos[8022]=25;
cos[8023]=25;
cos[8024]=25;
cos[8025]=25;
cos[8026]=25;
cos[8027]=25;
cos[8028]=25;
cos[8029]=25;
cos[8030]=26;
cos[8031]=26;
cos[8032]=26;
cos[8033]=26;
cos[8034]=26;
cos[8035]=26;
cos[8036]=26;
cos[8037]=26;
cos[8038]=26;
cos[8039]=26;
cos[8040]=26;
cos[8041]=26;
cos[8042]=26;
cos[8043]=26;
cos[8044]=26;
cos[8045]=26;
cos[8046]=26;
cos[8047]=26;
cos[8048]=26;
cos[8049]=26;
cos[8050]=26;
cos[8051]=27;
cos[8052]=27;
cos[8053]=27;
cos[8054]=27;
cos[8055]=27;
cos[8056]=27;
cos[8057]=27;
cos[8058]=27;
cos[8059]=27;
cos[8060]=27;
cos[8061]=27;
cos[8062]=27;
cos[8063]=27;
cos[8064]=27;
cos[8065]=27;
cos[8066]=27;
cos[8067]=27;
cos[8068]=27;
cos[8069]=27;
cos[8070]=27;
cos[8071]=27;
cos[8072]=27;
cos[8073]=28;
cos[8074]=28;
cos[8075]=28;
cos[8076]=28;
cos[8077]=28;
cos[8078]=28;
cos[8079]=28;
cos[8080]=28;
cos[8081]=28;
cos[8082]=28;
cos[8083]=28;
cos[8084]=28;
cos[8085]=28;
cos[8086]=28;
cos[8087]=28;
cos[8088]=28;
cos[8089]=28;
cos[8090]=28;
cos[8091]=28;
cos[8092]=28;
cos[8093]=28;
cos[8094]=28;
cos[8095]=29;
cos[8096]=29;
cos[8097]=29;
cos[8098]=29;
cos[8099]=29;
cos[8100]=29;
cos[8101]=29;
cos[8102]=29;
cos[8103]=29;
cos[8104]=29;
cos[8105]=29;
cos[8106]=29;
cos[8107]=29;
cos[8108]=29;
cos[8109]=29;
cos[8110]=29;
cos[8111]=29;
cos[8112]=29;
cos[8113]=29;
cos[8114]=29;
cos[8115]=29;
cos[8116]=29;
cos[8117]=30;
cos[8118]=30;
cos[8119]=30;
cos[8120]=30;
cos[8121]=30;
cos[8122]=30;
cos[8123]=30;
cos[8124]=30;
cos[8125]=30;
cos[8126]=30;
cos[8127]=30;
cos[8128]=30;
cos[8129]=30;
cos[8130]=30;
cos[8131]=30;
cos[8132]=30;
cos[8133]=30;
cos[8134]=30;
cos[8135]=30;
cos[8136]=30;
cos[8137]=30;
cos[8138]=30;
cos[8139]=31;
cos[8140]=31;
cos[8141]=31;
cos[8142]=31;
cos[8143]=31;
cos[8144]=31;
cos[8145]=31;
cos[8146]=31;
cos[8147]=31;
cos[8148]=31;
cos[8149]=31;
cos[8150]=31;
cos[8151]=31;
cos[8152]=31;
cos[8153]=31;
cos[8154]=31;
cos[8155]=31;
cos[8156]=31;
cos[8157]=31;
cos[8158]=31;
cos[8159]=31;
cos[8160]=31;
cos[8161]=32;
cos[8162]=32;
cos[8163]=32;
cos[8164]=32;
cos[8165]=32;
cos[8166]=32;
cos[8167]=32;
cos[8168]=32;
cos[8169]=32;
cos[8170]=32;
cos[8171]=32;
cos[8172]=32;
cos[8173]=32;
cos[8174]=32;
cos[8175]=32;
cos[8176]=32;
cos[8177]=32;
cos[8178]=32;
cos[8179]=32;
cos[8180]=32;
cos[8181]=32;
cos[8182]=32;
cos[8183]=33;
cos[8184]=33;
cos[8185]=33;
cos[8186]=33;
cos[8187]=33;
cos[8188]=33;
cos[8189]=33;
cos[8190]=33;
cos[8191]=33;
cos[8192]=33;
cos[8193]=33;
cos[8194]=33;
cos[8195]=33;
cos[8196]=33;
cos[8197]=33;
cos[8198]=33;
cos[8199]=33;
cos[8200]=33;
cos[8201]=33;
cos[8202]=33;
cos[8203]=33;
cos[8204]=33;
cos[8205]=33;
cos[8206]=34;
cos[8207]=34;
cos[8208]=34;
cos[8209]=34;
cos[8210]=34;
cos[8211]=34;
cos[8212]=34;
cos[8213]=34;
cos[8214]=34;
cos[8215]=34;
cos[8216]=34;
cos[8217]=34;
cos[8218]=34;
cos[8219]=34;
cos[8220]=34;
cos[8221]=34;
cos[8222]=34;
cos[8223]=34;
cos[8224]=34;
cos[8225]=34;
cos[8226]=34;
cos[8227]=34;
cos[8228]=35;
cos[8229]=35;
cos[8230]=35;
cos[8231]=35;
cos[8232]=35;
cos[8233]=35;
cos[8234]=35;
cos[8235]=35;
cos[8236]=35;
cos[8237]=35;
cos[8238]=35;
cos[8239]=35;
cos[8240]=35;
cos[8241]=35;
cos[8242]=35;
cos[8243]=35;
cos[8244]=35;
cos[8245]=35;
cos[8246]=35;
cos[8247]=35;
cos[8248]=35;
cos[8249]=35;
cos[8250]=35;
cos[8251]=36;
cos[8252]=36;
cos[8253]=36;
cos[8254]=36;
cos[8255]=36;
cos[8256]=36;
cos[8257]=36;
cos[8258]=36;
cos[8259]=36;
cos[8260]=36;
cos[8261]=36;
cos[8262]=36;
cos[8263]=36;
cos[8264]=36;
cos[8265]=36;
cos[8266]=36;
cos[8267]=36;
cos[8268]=36;
cos[8269]=36;
cos[8270]=36;
cos[8271]=36;
cos[8272]=36;
cos[8273]=36;
cos[8274]=37;
cos[8275]=37;
cos[8276]=37;
cos[8277]=37;
cos[8278]=37;
cos[8279]=37;
cos[8280]=37;
cos[8281]=37;
cos[8282]=37;
cos[8283]=37;
cos[8284]=37;
cos[8285]=37;
cos[8286]=37;
cos[8287]=37;
cos[8288]=37;
cos[8289]=37;
cos[8290]=37;
cos[8291]=37;
cos[8292]=37;
cos[8293]=37;
cos[8294]=37;
cos[8295]=37;
cos[8296]=37;
cos[8297]=38;
cos[8298]=38;
cos[8299]=38;
cos[8300]=38;
cos[8301]=38;
cos[8302]=38;
cos[8303]=38;
cos[8304]=38;
cos[8305]=38;
cos[8306]=38;
cos[8307]=38;
cos[8308]=38;
cos[8309]=38;
cos[8310]=38;
cos[8311]=38;
cos[8312]=38;
cos[8313]=38;
cos[8314]=38;
cos[8315]=38;
cos[8316]=38;
cos[8317]=38;
cos[8318]=38;
cos[8319]=38;
cos[8320]=38;
cos[8321]=39;
cos[8322]=39;
cos[8323]=39;
cos[8324]=39;
cos[8325]=39;
cos[8326]=39;
cos[8327]=39;
cos[8328]=39;
cos[8329]=39;
cos[8330]=39;
cos[8331]=39;
cos[8332]=39;
cos[8333]=39;
cos[8334]=39;
cos[8335]=39;
cos[8336]=39;
cos[8337]=39;
cos[8338]=39;
cos[8339]=39;
cos[8340]=39;
cos[8341]=39;
cos[8342]=39;
cos[8343]=39;
cos[8344]=40;
cos[8345]=40;
cos[8346]=40;
cos[8347]=40;
cos[8348]=40;
cos[8349]=40;
cos[8350]=40;
cos[8351]=40;
cos[8352]=40;
cos[8353]=40;
cos[8354]=40;
cos[8355]=40;
cos[8356]=40;
cos[8357]=40;
cos[8358]=40;
cos[8359]=40;
cos[8360]=40;
cos[8361]=40;
cos[8362]=40;
cos[8363]=40;
cos[8364]=40;
cos[8365]=40;
cos[8366]=40;
cos[8367]=40;
cos[8368]=41;
cos[8369]=41;
cos[8370]=41;
cos[8371]=41;
cos[8372]=41;
cos[8373]=41;
cos[8374]=41;
cos[8375]=41;
cos[8376]=41;
cos[8377]=41;
cos[8378]=41;
cos[8379]=41;
cos[8380]=41;
cos[8381]=41;
cos[8382]=41;
cos[8383]=41;
cos[8384]=41;
cos[8385]=41;
cos[8386]=41;
cos[8387]=41;
cos[8388]=41;
cos[8389]=41;
cos[8390]=41;
cos[8391]=41;
cos[8392]=42;
cos[8393]=42;
cos[8394]=42;
cos[8395]=42;
cos[8396]=42;
cos[8397]=42;
cos[8398]=42;
cos[8399]=42;
cos[8400]=42;
cos[8401]=42;
cos[8402]=42;
cos[8403]=42;
cos[8404]=42;
cos[8405]=42;
cos[8406]=42;
cos[8407]=42;
cos[8408]=42;
cos[8409]=42;
cos[8410]=42;
cos[8411]=42;
cos[8412]=42;
cos[8413]=42;
cos[8414]=42;
cos[8415]=42;
cos[8416]=43;
cos[8417]=43;
cos[8418]=43;
cos[8419]=43;
cos[8420]=43;
cos[8421]=43;
cos[8422]=43;
cos[8423]=43;
cos[8424]=43;
cos[8425]=43;
cos[8426]=43;
cos[8427]=43;
cos[8428]=43;
cos[8429]=43;
cos[8430]=43;
cos[8431]=43;
cos[8432]=43;
cos[8433]=43;
cos[8434]=43;
cos[8435]=43;
cos[8436]=43;
cos[8437]=43;
cos[8438]=43;
cos[8439]=43;
cos[8440]=44;
cos[8441]=44;
cos[8442]=44;
cos[8443]=44;
cos[8444]=44;
cos[8445]=44;
cos[8446]=44;
cos[8447]=44;
cos[8448]=44;
cos[8449]=44;
cos[8450]=44;
cos[8451]=44;
cos[8452]=44;
cos[8453]=44;
cos[8454]=44;
cos[8455]=44;
cos[8456]=44;
cos[8457]=44;
cos[8458]=44;
cos[8459]=44;
cos[8460]=44;
cos[8461]=44;
cos[8462]=44;
cos[8463]=44;
cos[8464]=44;
cos[8465]=45;
cos[8466]=45;
cos[8467]=45;
cos[8468]=45;
cos[8469]=45;
cos[8470]=45;
cos[8471]=45;
cos[8472]=45;
cos[8473]=45;
cos[8474]=45;
cos[8475]=45;
cos[8476]=45;
cos[8477]=45;
cos[8478]=45;
cos[8479]=45;
cos[8480]=45;
cos[8481]=45;
cos[8482]=45;
cos[8483]=45;
cos[8484]=45;
cos[8485]=45;
cos[8486]=45;
cos[8487]=45;
cos[8488]=45;
cos[8489]=45;
cos[8490]=46;
cos[8491]=46;
cos[8492]=46;
cos[8493]=46;
cos[8494]=46;
cos[8495]=46;
cos[8496]=46;
cos[8497]=46;
cos[8498]=46;
cos[8499]=46;
cos[8500]=46;
cos[8501]=46;
cos[8502]=46;
cos[8503]=46;
cos[8504]=46;
cos[8505]=46;
cos[8506]=46;
cos[8507]=46;
cos[8508]=46;
cos[8509]=46;
cos[8510]=46;
cos[8511]=46;
cos[8512]=46;
cos[8513]=46;
cos[8514]=46;
cos[8515]=47;
cos[8516]=47;
cos[8517]=47;
cos[8518]=47;
cos[8519]=47;
cos[8520]=47;
cos[8521]=47;
cos[8522]=47;
cos[8523]=47;
cos[8524]=47;
cos[8525]=47;
cos[8526]=47;
cos[8527]=47;
cos[8528]=47;
cos[8529]=47;
cos[8530]=47;
cos[8531]=47;
cos[8532]=47;
cos[8533]=47;
cos[8534]=47;
cos[8535]=47;
cos[8536]=47;
cos[8537]=47;
cos[8538]=47;
cos[8539]=47;
cos[8540]=47;
cos[8541]=48;
cos[8542]=48;
cos[8543]=48;
cos[8544]=48;
cos[8545]=48;
cos[8546]=48;
cos[8547]=48;
cos[8548]=48;
cos[8549]=48;
cos[8550]=48;
cos[8551]=48;
cos[8552]=48;
cos[8553]=48;
cos[8554]=48;
cos[8555]=48;
cos[8556]=48;
cos[8557]=48;
cos[8558]=48;
cos[8559]=48;
cos[8560]=48;
cos[8561]=48;
cos[8562]=48;
cos[8563]=48;
cos[8564]=48;
cos[8565]=48;
cos[8566]=49;
cos[8567]=49;
cos[8568]=49;
cos[8569]=49;
cos[8570]=49;
cos[8571]=49;
cos[8572]=49;
cos[8573]=49;
cos[8574]=49;
cos[8575]=49;
cos[8576]=49;
cos[8577]=49;
cos[8578]=49;
cos[8579]=49;
cos[8580]=49;
cos[8581]=49;
cos[8582]=49;
cos[8583]=49;
cos[8584]=49;
cos[8585]=49;
cos[8586]=49;
cos[8587]=49;
cos[8588]=49;
cos[8589]=49;
cos[8590]=49;
cos[8591]=49;
cos[8592]=49;
cos[8593]=50;
cos[8594]=50;
cos[8595]=50;
cos[8596]=50;
cos[8597]=50;
cos[8598]=50;
cos[8599]=50;
cos[8600]=50;
cos[8601]=50;
cos[8602]=50;
cos[8603]=50;
cos[8604]=50;
cos[8605]=50;
cos[8606]=50;
cos[8607]=50;
cos[8608]=50;
cos[8609]=50;
cos[8610]=50;
cos[8611]=50;
cos[8612]=50;
cos[8613]=50;
cos[8614]=50;
cos[8615]=50;
cos[8616]=50;
cos[8617]=50;
cos[8618]=50;
cos[8619]=51;
cos[8620]=51;
cos[8621]=51;
cos[8622]=51;
cos[8623]=51;
cos[8624]=51;
cos[8625]=51;
cos[8626]=51;
cos[8627]=51;
cos[8628]=51;
cos[8629]=51;
cos[8630]=51;
cos[8631]=51;
cos[8632]=51;
cos[8633]=51;
cos[8634]=51;
cos[8635]=51;
cos[8636]=51;
cos[8637]=51;
cos[8638]=51;
cos[8639]=51;
cos[8640]=51;
cos[8641]=51;
cos[8642]=51;
cos[8643]=51;
cos[8644]=51;
cos[8645]=51;
cos[8646]=52;
cos[8647]=52;
cos[8648]=52;
cos[8649]=52;
cos[8650]=52;
cos[8651]=52;
cos[8652]=52;
cos[8653]=52;
cos[8654]=52;
cos[8655]=52;
cos[8656]=52;
cos[8657]=52;
cos[8658]=52;
cos[8659]=52;
cos[8660]=52;
cos[8661]=52;
cos[8662]=52;
cos[8663]=52;
cos[8664]=52;
cos[8665]=52;
cos[8666]=52;
cos[8667]=52;
cos[8668]=52;
cos[8669]=52;
cos[8670]=52;
cos[8671]=52;
cos[8672]=52;
cos[8673]=53;
cos[8674]=53;
cos[8675]=53;
cos[8676]=53;
cos[8677]=53;
cos[8678]=53;
cos[8679]=53;
cos[8680]=53;
cos[8681]=53;
cos[8682]=53;
cos[8683]=53;
cos[8684]=53;
cos[8685]=53;
cos[8686]=53;
cos[8687]=53;
cos[8688]=53;
cos[8689]=53;
cos[8690]=53;
cos[8691]=53;
cos[8692]=53;
cos[8693]=53;
cos[8694]=53;
cos[8695]=53;
cos[8696]=53;
cos[8697]=53;
cos[8698]=53;
cos[8699]=53;
cos[8700]=53;
cos[8701]=54;
cos[8702]=54;
cos[8703]=54;
cos[8704]=54;
cos[8705]=54;
cos[8706]=54;
cos[8707]=54;
cos[8708]=54;
cos[8709]=54;
cos[8710]=54;
cos[8711]=54;
cos[8712]=54;
cos[8713]=54;
cos[8714]=54;
cos[8715]=54;
cos[8716]=54;
cos[8717]=54;
cos[8718]=54;
cos[8719]=54;
cos[8720]=54;
cos[8721]=54;
cos[8722]=54;
cos[8723]=54;
cos[8724]=54;
cos[8725]=54;
cos[8726]=54;
cos[8727]=54;
cos[8728]=54;
cos[8729]=55;
cos[8730]=55;
cos[8731]=55;
cos[8732]=55;
cos[8733]=55;
cos[8734]=55;
cos[8735]=55;
cos[8736]=55;
cos[8737]=55;
cos[8738]=55;
cos[8739]=55;
cos[8740]=55;
cos[8741]=55;
cos[8742]=55;
cos[8743]=55;
cos[8744]=55;
cos[8745]=55;
cos[8746]=55;
cos[8747]=55;
cos[8748]=55;
cos[8749]=55;
cos[8750]=55;
cos[8751]=55;
cos[8752]=55;
cos[8753]=55;
cos[8754]=55;
cos[8755]=55;
cos[8756]=55;
cos[8757]=55;
cos[8758]=56;
cos[8759]=56;
cos[8760]=56;
cos[8761]=56;
cos[8762]=56;
cos[8763]=56;
cos[8764]=56;
cos[8765]=56;
cos[8766]=56;
cos[8767]=56;
cos[8768]=56;
cos[8769]=56;
cos[8770]=56;
cos[8771]=56;
cos[8772]=56;
cos[8773]=56;
cos[8774]=56;
cos[8775]=56;
cos[8776]=56;
cos[8777]=56;
cos[8778]=56;
cos[8779]=56;
cos[8780]=56;
cos[8781]=56;
cos[8782]=56;
cos[8783]=56;
cos[8784]=56;
cos[8785]=56;
cos[8786]=56;
cos[8787]=57;
cos[8788]=57;
cos[8789]=57;
cos[8790]=57;
cos[8791]=57;
cos[8792]=57;
cos[8793]=57;
cos[8794]=57;
cos[8795]=57;
cos[8796]=57;
cos[8797]=57;
cos[8798]=57;
cos[8799]=57;
cos[8800]=57;
cos[8801]=57;
cos[8802]=57;
cos[8803]=57;
cos[8804]=57;
cos[8805]=57;
cos[8806]=57;
cos[8807]=57;
cos[8808]=57;
cos[8809]=57;
cos[8810]=57;
cos[8811]=57;
cos[8812]=57;
cos[8813]=57;
cos[8814]=57;
cos[8815]=57;
cos[8816]=57;
cos[8817]=58;
cos[8818]=58;
cos[8819]=58;
cos[8820]=58;
cos[8821]=58;
cos[8822]=58;
cos[8823]=58;
cos[8824]=58;
cos[8825]=58;
cos[8826]=58;
cos[8827]=58;
cos[8828]=58;
cos[8829]=58;
cos[8830]=58;
cos[8831]=58;
cos[8832]=58;
cos[8833]=58;
cos[8834]=58;
cos[8835]=58;
cos[8836]=58;
cos[8837]=58;
cos[8838]=58;
cos[8839]=58;
cos[8840]=58;
cos[8841]=58;
cos[8842]=58;
cos[8843]=58;
cos[8844]=58;
cos[8845]=58;
cos[8846]=58;
cos[8847]=59;
cos[8848]=59;
cos[8849]=59;
cos[8850]=59;
cos[8851]=59;
cos[8852]=59;
cos[8853]=59;
cos[8854]=59;
cos[8855]=59;
cos[8856]=59;
cos[8857]=59;
cos[8858]=59;
cos[8859]=59;
cos[8860]=59;
cos[8861]=59;
cos[8862]=59;
cos[8863]=59;
cos[8864]=59;
cos[8865]=59;
cos[8866]=59;
cos[8867]=59;
cos[8868]=59;
cos[8869]=59;
cos[8870]=59;
cos[8871]=59;
cos[8872]=59;
cos[8873]=59;
cos[8874]=59;
cos[8875]=59;
cos[8876]=59;
cos[8877]=59;
cos[8878]=60;
cos[8879]=60;
cos[8880]=60;
cos[8881]=60;
cos[8882]=60;
cos[8883]=60;
cos[8884]=60;
cos[8885]=60;
cos[8886]=60;
cos[8887]=60;
cos[8888]=60;
cos[8889]=60;
cos[8890]=60;
cos[8891]=60;
cos[8892]=60;
cos[8893]=60;
cos[8894]=60;
cos[8895]=60;
cos[8896]=60;
cos[8897]=60;
cos[8898]=60;
cos[8899]=60;
cos[8900]=60;
cos[8901]=60;
cos[8902]=60;
cos[8903]=60;
cos[8904]=60;
cos[8905]=60;
cos[8906]=60;
cos[8907]=60;
cos[8908]=60;
cos[8909]=60;
cos[8910]=61;
cos[8911]=61;
cos[8912]=61;
cos[8913]=61;
cos[8914]=61;
cos[8915]=61;
cos[8916]=61;
cos[8917]=61;
cos[8918]=61;
cos[8919]=61;
cos[8920]=61;
cos[8921]=61;
cos[8922]=61;
cos[8923]=61;
cos[8924]=61;
cos[8925]=61;
cos[8926]=61;
cos[8927]=61;
cos[8928]=61;
cos[8929]=61;
cos[8930]=61;
cos[8931]=61;
cos[8932]=61;
cos[8933]=61;
cos[8934]=61;
cos[8935]=61;
cos[8936]=61;
cos[8937]=61;
cos[8938]=61;
cos[8939]=61;
cos[8940]=61;
cos[8941]=61;
cos[8942]=61;
cos[8943]=62;
cos[8944]=62;
cos[8945]=62;
cos[8946]=62;
cos[8947]=62;
cos[8948]=62;
cos[8949]=62;
cos[8950]=62;
cos[8951]=62;
cos[8952]=62;
cos[8953]=62;
cos[8954]=62;
cos[8955]=62;
cos[8956]=62;
cos[8957]=62;
cos[8958]=62;
cos[8959]=62;
cos[8960]=62;
cos[8961]=62;
cos[8962]=62;
cos[8963]=62;
cos[8964]=62;
cos[8965]=62;
cos[8966]=62;
cos[8967]=62;
cos[8968]=62;
cos[8969]=62;
cos[8970]=62;
cos[8971]=62;
cos[8972]=62;
cos[8973]=62;
cos[8974]=62;
cos[8975]=62;
cos[8976]=63;
cos[8977]=63;
cos[8978]=63;
cos[8979]=63;
cos[8980]=63;
cos[8981]=63;
cos[8982]=63;
cos[8983]=63;
cos[8984]=63;
cos[8985]=63;
cos[8986]=63;
cos[8987]=63;
cos[8988]=63;
cos[8989]=63;
cos[8990]=63;
cos[8991]=63;
cos[8992]=63;
cos[8993]=63;
cos[8994]=63;
cos[8995]=63;
cos[8996]=63;
cos[8997]=63;
cos[8998]=63;
cos[8999]=63;
cos[9000]=63;
cos[9001]=63;
cos[9002]=63;
cos[9003]=63;
cos[9004]=63;
cos[9005]=63;
cos[9006]=63;
cos[9007]=63;
cos[9008]=63;
cos[9009]=63;
cos[9010]=63;
cos[9011]=64;
cos[9012]=64;
cos[9013]=64;
cos[9014]=64;
cos[9015]=64;
cos[9016]=64;
cos[9017]=64;
cos[9018]=64;
cos[9019]=64;
cos[9020]=64;
cos[9021]=64;
cos[9022]=64;
cos[9023]=64;
cos[9024]=64;
cos[9025]=64;
cos[9026]=64;
cos[9027]=64;
cos[9028]=64;
cos[9029]=64;
cos[9030]=64;
cos[9031]=64;
cos[9032]=64;
cos[9033]=64;
cos[9034]=64;
cos[9035]=64;
cos[9036]=64;
cos[9037]=64;
cos[9038]=64;
cos[9039]=64;
cos[9040]=64;
cos[9041]=64;
cos[9042]=64;
cos[9043]=64;
cos[9044]=64;
cos[9045]=64;
cos[9046]=65;
cos[9047]=65;
cos[9048]=65;
cos[9049]=65;
cos[9050]=65;
cos[9051]=65;
cos[9052]=65;
cos[9053]=65;
cos[9054]=65;
cos[9055]=65;
cos[9056]=65;
cos[9057]=65;
cos[9058]=65;
cos[9059]=65;
cos[9060]=65;
cos[9061]=65;
cos[9062]=65;
cos[9063]=65;
cos[9064]=65;
cos[9065]=65;
cos[9066]=65;
cos[9067]=65;
cos[9068]=65;
cos[9069]=65;
cos[9070]=65;
cos[9071]=65;
cos[9072]=65;
cos[9073]=65;
cos[9074]=65;
cos[9075]=65;
cos[9076]=65;
cos[9077]=65;
cos[9078]=65;
cos[9079]=65;
cos[9080]=65;
cos[9081]=65;
cos[9082]=65;
cos[9083]=66;
cos[9084]=66;
cos[9085]=66;
cos[9086]=66;
cos[9087]=66;
cos[9088]=66;
cos[9089]=66;
cos[9090]=66;
cos[9091]=66;
cos[9092]=66;
cos[9093]=66;
cos[9094]=66;
cos[9095]=66;
cos[9096]=66;
cos[9097]=66;
cos[9098]=66;
cos[9099]=66;
cos[9100]=66;
cos[9101]=66;
cos[9102]=66;
cos[9103]=66;
cos[9104]=66;
cos[9105]=66;
cos[9106]=66;
cos[9107]=66;
cos[9108]=66;
cos[9109]=66;
cos[9110]=66;
cos[9111]=66;
cos[9112]=66;
cos[9113]=66;
cos[9114]=66;
cos[9115]=66;
cos[9116]=66;
cos[9117]=66;
cos[9118]=66;
cos[9119]=66;
cos[9120]=66;
cos[9121]=67;
cos[9122]=67;
cos[9123]=67;
cos[9124]=67;
cos[9125]=67;
cos[9126]=67;
cos[9127]=67;
cos[9128]=67;
cos[9129]=67;
cos[9130]=67;
cos[9131]=67;
cos[9132]=67;
cos[9133]=67;
cos[9134]=67;
cos[9135]=67;
cos[9136]=67;
cos[9137]=67;
cos[9138]=67;
cos[9139]=67;
cos[9140]=67;
cos[9141]=67;
cos[9142]=67;
cos[9143]=67;
cos[9144]=67;
cos[9145]=67;
cos[9146]=67;
cos[9147]=67;
cos[9148]=67;
cos[9149]=67;
cos[9150]=67;
cos[9151]=67;
cos[9152]=67;
cos[9153]=67;
cos[9154]=67;
cos[9155]=67;
cos[9156]=67;
cos[9157]=67;
cos[9158]=67;
cos[9159]=67;
cos[9160]=67;
cos[9161]=68;
cos[9162]=68;
cos[9163]=68;
cos[9164]=68;
cos[9165]=68;
cos[9166]=68;
cos[9167]=68;
cos[9168]=68;
cos[9169]=68;
cos[9170]=68;
cos[9171]=68;
cos[9172]=68;
cos[9173]=68;
cos[9174]=68;
cos[9175]=68;
cos[9176]=68;
cos[9177]=68;
cos[9178]=68;
cos[9179]=68;
cos[9180]=68;
cos[9181]=68;
cos[9182]=68;
cos[9183]=68;
cos[9184]=68;
cos[9185]=68;
cos[9186]=68;
cos[9187]=68;
cos[9188]=68;
cos[9189]=68;
cos[9190]=68;
cos[9191]=68;
cos[9192]=68;
cos[9193]=68;
cos[9194]=68;
cos[9195]=68;
cos[9196]=68;
cos[9197]=68;
cos[9198]=68;
cos[9199]=68;
cos[9200]=68;
cos[9201]=68;
cos[9202]=69;
cos[9203]=69;
cos[9204]=69;
cos[9205]=69;
cos[9206]=69;
cos[9207]=69;
cos[9208]=69;
cos[9209]=69;
cos[9210]=69;
cos[9211]=69;
cos[9212]=69;
cos[9213]=69;
cos[9214]=69;
cos[9215]=69;
cos[9216]=69;
cos[9217]=69;
cos[9218]=69;
cos[9219]=69;
cos[9220]=69;
cos[9221]=69;
cos[9222]=69;
cos[9223]=69;
cos[9224]=69;
cos[9225]=69;
cos[9226]=69;
cos[9227]=69;
cos[9228]=69;
cos[9229]=69;
cos[9230]=69;
cos[9231]=69;
cos[9232]=69;
cos[9233]=69;
cos[9234]=69;
cos[9235]=69;
cos[9236]=69;
cos[9237]=69;
cos[9238]=69;
cos[9239]=69;
cos[9240]=69;
cos[9241]=69;
cos[9242]=69;
cos[9243]=69;
cos[9244]=69;
cos[9245]=69;
cos[9246]=70;
cos[9247]=70;
cos[9248]=70;
cos[9249]=70;
cos[9250]=70;
cos[9251]=70;
cos[9252]=70;
cos[9253]=70;
cos[9254]=70;
cos[9255]=70;
cos[9256]=70;
cos[9257]=70;
cos[9258]=70;
cos[9259]=70;
cos[9260]=70;
cos[9261]=70;
cos[9262]=70;
cos[9263]=70;
cos[9264]=70;
cos[9265]=70;
cos[9266]=70;
cos[9267]=70;
cos[9268]=70;
cos[9269]=70;
cos[9270]=70;
cos[9271]=70;
cos[9272]=70;
cos[9273]=70;
cos[9274]=70;
cos[9275]=70;
cos[9276]=70;
cos[9277]=70;
cos[9278]=70;
cos[9279]=70;
cos[9280]=70;
cos[9281]=70;
cos[9282]=70;
cos[9283]=70;
cos[9284]=70;
cos[9285]=70;
cos[9286]=70;
cos[9287]=70;
cos[9288]=70;
cos[9289]=70;
cos[9290]=70;
cos[9291]=71;
cos[9292]=71;
cos[9293]=71;
cos[9294]=71;
cos[9295]=71;
cos[9296]=71;
cos[9297]=71;
cos[9298]=71;
cos[9299]=71;
cos[9300]=71;
cos[9301]=71;
cos[9302]=71;
cos[9303]=71;
cos[9304]=71;
cos[9305]=71;
cos[9306]=71;
cos[9307]=71;
cos[9308]=71;
cos[9309]=71;
cos[9310]=71;
cos[9311]=71;
cos[9312]=71;
cos[9313]=71;
cos[9314]=71;
cos[9315]=71;
cos[9316]=71;
cos[9317]=71;
cos[9318]=71;
cos[9319]=71;
cos[9320]=71;
cos[9321]=71;
cos[9322]=71;
cos[9323]=71;
cos[9324]=71;
cos[9325]=71;
cos[9326]=71;
cos[9327]=71;
cos[9328]=71;
cos[9329]=71;
cos[9330]=71;
cos[9331]=71;
cos[9332]=71;
cos[9333]=71;
cos[9334]=71;
cos[9335]=71;
cos[9336]=71;
cos[9337]=71;
cos[9338]=71;
cos[9339]=71;
cos[9340]=72;
cos[9341]=72;
cos[9342]=72;
cos[9343]=72;
cos[9344]=72;
cos[9345]=72;
cos[9346]=72;
cos[9347]=72;
cos[9348]=72;
cos[9349]=72;
cos[9350]=72;
cos[9351]=72;
cos[9352]=72;
cos[9353]=72;
cos[9354]=72;
cos[9355]=72;
cos[9356]=72;
cos[9357]=72;
cos[9358]=72;
cos[9359]=72;
cos[9360]=72;
cos[9361]=72;
cos[9362]=72;
cos[9363]=72;
cos[9364]=72;
cos[9365]=72;
cos[9366]=72;
cos[9367]=72;
cos[9368]=72;
cos[9369]=72;
cos[9370]=72;
cos[9371]=72;
cos[9372]=72;
cos[9373]=72;
cos[9374]=72;
cos[9375]=72;
cos[9376]=72;
cos[9377]=72;
cos[9378]=72;
cos[9379]=72;
cos[9380]=72;
cos[9381]=72;
cos[9382]=72;
cos[9383]=72;
cos[9384]=72;
cos[9385]=72;
cos[9386]=72;
cos[9387]=72;
cos[9388]=72;
cos[9389]=72;
cos[9390]=72;
cos[9391]=72;
cos[9392]=72;
cos[9393]=73;
cos[9394]=73;
cos[9395]=73;
cos[9396]=73;
cos[9397]=73;
cos[9398]=73;
cos[9399]=73;
cos[9400]=73;
cos[9401]=73;
cos[9402]=73;
cos[9403]=73;
cos[9404]=73;
cos[9405]=73;
cos[9406]=73;
cos[9407]=73;
cos[9408]=73;
cos[9409]=73;
cos[9410]=73;
cos[9411]=73;
cos[9412]=73;
cos[9413]=73;
cos[9414]=73;
cos[9415]=73;
cos[9416]=73;
cos[9417]=73;
cos[9418]=73;
cos[9419]=73;
cos[9420]=73;
cos[9421]=73;
cos[9422]=73;
cos[9423]=73;
cos[9424]=73;
cos[9425]=73;
cos[9426]=73;
cos[9427]=73;
cos[9428]=73;
cos[9429]=73;
cos[9430]=73;
cos[9431]=73;
cos[9432]=73;
cos[9433]=73;
cos[9434]=73;
cos[9435]=73;
cos[9436]=73;
cos[9437]=73;
cos[9438]=73;
cos[9439]=73;
cos[9440]=73;
cos[9441]=73;
cos[9442]=73;
cos[9443]=73;
cos[9444]=73;
cos[9445]=73;
cos[9446]=73;
cos[9447]=73;
cos[9448]=73;
cos[9449]=73;
cos[9450]=74;
cos[9451]=74;
cos[9452]=74;
cos[9453]=74;
cos[9454]=74;
cos[9455]=74;
cos[9456]=74;
cos[9457]=74;
cos[9458]=74;
cos[9459]=74;
cos[9460]=74;
cos[9461]=74;
cos[9462]=74;
cos[9463]=74;
cos[9464]=74;
cos[9465]=74;
cos[9466]=74;
cos[9467]=74;
cos[9468]=74;
cos[9469]=74;
cos[9470]=74;
cos[9471]=74;
cos[9472]=74;
cos[9473]=74;
cos[9474]=74;
cos[9475]=74;
cos[9476]=74;
cos[9477]=74;
cos[9478]=74;
cos[9479]=74;
cos[9480]=74;
cos[9481]=74;
cos[9482]=74;
cos[9483]=74;
cos[9484]=74;
cos[9485]=74;
cos[9486]=74;
cos[9487]=74;
cos[9488]=74;
cos[9489]=74;
cos[9490]=74;
cos[9491]=74;
cos[9492]=74;
cos[9493]=74;
cos[9494]=74;
cos[9495]=74;
cos[9496]=74;
cos[9497]=74;
cos[9498]=74;
cos[9499]=74;
cos[9500]=74;
cos[9501]=74;
cos[9502]=74;
cos[9503]=74;
cos[9504]=74;
cos[9505]=74;
cos[9506]=74;
cos[9507]=74;
cos[9508]=74;
cos[9509]=74;
cos[9510]=74;
cos[9511]=74;
cos[9512]=74;
cos[9513]=74;
cos[9514]=75;
cos[9515]=75;
cos[9516]=75;
cos[9517]=75;
cos[9518]=75;
cos[9519]=75;
cos[9520]=75;
cos[9521]=75;
cos[9522]=75;
cos[9523]=75;
cos[9524]=75;
cos[9525]=75;
cos[9526]=75;
cos[9527]=75;
cos[9528]=75;
cos[9529]=75;
cos[9530]=75;
cos[9531]=75;
cos[9532]=75;
cos[9533]=75;
cos[9534]=75;
cos[9535]=75;
cos[9536]=75;
cos[9537]=75;
cos[9538]=75;
cos[9539]=75;
cos[9540]=75;
cos[9541]=75;
cos[9542]=75;
cos[9543]=75;
cos[9544]=75;
cos[9545]=75;
cos[9546]=75;
cos[9547]=75;
cos[9548]=75;
cos[9549]=75;
cos[9550]=75;
cos[9551]=75;
cos[9552]=75;
cos[9553]=75;
cos[9554]=75;
cos[9555]=75;
cos[9556]=75;
cos[9557]=75;
cos[9558]=75;
cos[9559]=75;
cos[9560]=75;
cos[9561]=75;
cos[9562]=75;
cos[9563]=75;
cos[9564]=75;
cos[9565]=75;
cos[9566]=75;
cos[9567]=75;
cos[9568]=75;
cos[9569]=75;
cos[9570]=75;
cos[9571]=75;
cos[9572]=75;
cos[9573]=75;
cos[9574]=75;
cos[9575]=75;
cos[9576]=75;
cos[9577]=75;
cos[9578]=75;
cos[9579]=75;
cos[9580]=75;
cos[9581]=75;
cos[9582]=75;
cos[9583]=75;
cos[9584]=75;
cos[9585]=75;
cos[9586]=75;
cos[9587]=76;
cos[9588]=76;
cos[9589]=76;
cos[9590]=76;
cos[9591]=76;
cos[9592]=76;
cos[9593]=76;
cos[9594]=76;
cos[9595]=76;
cos[9596]=76;
cos[9597]=76;
cos[9598]=76;
cos[9599]=76;
cos[9600]=76;
cos[9601]=76;
cos[9602]=76;
cos[9603]=76;
cos[9604]=76;
cos[9605]=76;
cos[9606]=76;
cos[9607]=76;
cos[9608]=76;
cos[9609]=76;
cos[9610]=76;
cos[9611]=76;
cos[9612]=76;
cos[9613]=76;
cos[9614]=76;
cos[9615]=76;
cos[9616]=76;
cos[9617]=76;
cos[9618]=76;
cos[9619]=76;
cos[9620]=76;
cos[9621]=76;
cos[9622]=76;
cos[9623]=76;
cos[9624]=76;
cos[9625]=76;
cos[9626]=76;
cos[9627]=76;
cos[9628]=76;
cos[9629]=76;
cos[9630]=76;
cos[9631]=76;
cos[9632]=76;
cos[9633]=76;
cos[9634]=76;
cos[9635]=76;
cos[9636]=76;
cos[9637]=76;
cos[9638]=76;
cos[9639]=76;
cos[9640]=76;
cos[9641]=76;
cos[9642]=76;
cos[9643]=76;
cos[9644]=76;
cos[9645]=76;
cos[9646]=76;
cos[9647]=76;
cos[9648]=76;
cos[9649]=76;
cos[9650]=76;
cos[9651]=76;
cos[9652]=76;
cos[9653]=76;
cos[9654]=76;
cos[9655]=76;
cos[9656]=76;
cos[9657]=76;
cos[9658]=76;
cos[9659]=76;
cos[9660]=76;
cos[9661]=76;
cos[9662]=76;
cos[9663]=76;
cos[9664]=76;
cos[9665]=76;
cos[9666]=76;
cos[9667]=76;
cos[9668]=76;
cos[9669]=76;
cos[9670]=76;
cos[9671]=76;
cos[9672]=76;
cos[9673]=76;
cos[9674]=76;
cos[9675]=77;
cos[9676]=77;
cos[9677]=77;
cos[9678]=77;
cos[9679]=77;
cos[9680]=77;
cos[9681]=77;
cos[9682]=77;
cos[9683]=77;
cos[9684]=77;
cos[9685]=77;
cos[9686]=77;
cos[9687]=77;
cos[9688]=77;
cos[9689]=77;
cos[9690]=77;
cos[9691]=77;
cos[9692]=77;
cos[9693]=77;
cos[9694]=77;
cos[9695]=77;
cos[9696]=77;
cos[9697]=77;
cos[9698]=77;
cos[9699]=77;
cos[9700]=77;
cos[9701]=77;
cos[9702]=77;
cos[9703]=77;
cos[9704]=77;
cos[9705]=77;
cos[9706]=77;
cos[9707]=77;
cos[9708]=77;
cos[9709]=77;
cos[9710]=77;
cos[9711]=77;
cos[9712]=77;
cos[9713]=77;
cos[9714]=77;
cos[9715]=77;
cos[9716]=77;
cos[9717]=77;
cos[9718]=77;
cos[9719]=77;
cos[9720]=77;
cos[9721]=77;
cos[9722]=77;
cos[9723]=77;
cos[9724]=77;
cos[9725]=77;
cos[9726]=77;
cos[9727]=77;
cos[9728]=77;
cos[9729]=77;
cos[9730]=77;
cos[9731]=77;
cos[9732]=77;
cos[9733]=77;
cos[9734]=77;
cos[9735]=77;
cos[9736]=77;
cos[9737]=77;
cos[9738]=77;
cos[9739]=77;
cos[9740]=77;
cos[9741]=77;
cos[9742]=77;
cos[9743]=77;
cos[9744]=77;
cos[9745]=77;
cos[9746]=77;
cos[9747]=77;
cos[9748]=77;
cos[9749]=77;
cos[9750]=77;
cos[9751]=77;
cos[9752]=77;
cos[9753]=77;
cos[9754]=77;
cos[9755]=77;
cos[9756]=77;
cos[9757]=77;
cos[9758]=77;
cos[9759]=77;
cos[9760]=77;
cos[9761]=77;
cos[9762]=77;
cos[9763]=77;
cos[9764]=77;
cos[9765]=77;
cos[9766]=77;
cos[9767]=77;
cos[9768]=77;
cos[9769]=77;
cos[9770]=77;
cos[9771]=77;
cos[9772]=77;
cos[9773]=77;
cos[9774]=77;
cos[9775]=77;
cos[9776]=77;
cos[9777]=77;
cos[9778]=77;
cos[9779]=77;
cos[9780]=77;
cos[9781]=77;
cos[9782]=77;
cos[9783]=77;
cos[9784]=77;
cos[9785]=77;
cos[9786]=77;
cos[9787]=77;
cos[9788]=77;
cos[9789]=77;
cos[9790]=77;
cos[9791]=77;
cos[9792]=77;
cos[9793]=77;
cos[9794]=77;
cos[9795]=77;
cos[9796]=77;
cos[9797]=77;
cos[9798]=77;
cos[9799]=78;
cos[9800]=78;
cos[9801]=78;
cos[9802]=78;
cos[9803]=78;
cos[9804]=78;
cos[9805]=78;
cos[9806]=78;
cos[9807]=78;
cos[9808]=78;
cos[9809]=78;
cos[9810]=78;
cos[9811]=78;
cos[9812]=78;
cos[9813]=78;
cos[9814]=78;
cos[9815]=78;
cos[9816]=78;
cos[9817]=78;
cos[9818]=78;
cos[9819]=78;
cos[9820]=78;
cos[9821]=78;
cos[9822]=78;
cos[9823]=78;
cos[9824]=78;
cos[9825]=78;
cos[9826]=78;
cos[9827]=78;
cos[9828]=78;
cos[9829]=78;
cos[9830]=78;
cos[9831]=78;
cos[9832]=78;
cos[9833]=78;
cos[9834]=78;
cos[9835]=78;
cos[9836]=78;
cos[9837]=78;
cos[9838]=78;
cos[9839]=78;
cos[9840]=78;
cos[9841]=78;
cos[9842]=78;
cos[9843]=78;
cos[9844]=78;
cos[9845]=78;
cos[9846]=78;
cos[9847]=78;
cos[9848]=78;
cos[9849]=78;
cos[9850]=78;
cos[9851]=78;
cos[9852]=78;
cos[9853]=78;
cos[9854]=78;
cos[9855]=78;
cos[9856]=78;
cos[9857]=78;
cos[9858]=78;
cos[9859]=78;
cos[9860]=78;
cos[9861]=78;
cos[9862]=78;
cos[9863]=78;
cos[9864]=78;
cos[9865]=78;
cos[9866]=78;
cos[9867]=78;
cos[9868]=78;
cos[9869]=78;
cos[9870]=78;
cos[9871]=78;
cos[9872]=78;
cos[9873]=78;
cos[9874]=78;
cos[9875]=78;
cos[9876]=78;
cos[9877]=78;
cos[9878]=78;
cos[9879]=78;
cos[9880]=78;
cos[9881]=78;
cos[9882]=78;
cos[9883]=78;
cos[9884]=78;
cos[9885]=78;
cos[9886]=78;
cos[9887]=78;
cos[9888]=78;
cos[9889]=78;
cos[9890]=78;
cos[9891]=78;
cos[9892]=78;
cos[9893]=78;
cos[9894]=78;
cos[9895]=78;
cos[9896]=78;
cos[9897]=78;
cos[9898]=78;
cos[9899]=78;
cos[9900]=78;
cos[9901]=78;
cos[9902]=78;
cos[9903]=78;
cos[9904]=78;
cos[9905]=78;
cos[9906]=78;
cos[9907]=78;
cos[9908]=78;
cos[9909]=78;
cos[9910]=78;
cos[9911]=78;
cos[9912]=78;
cos[9913]=78;
cos[9914]=78;
cos[9915]=78;
cos[9916]=78;
cos[9917]=78;
cos[9918]=78;
cos[9919]=78;
cos[9920]=78;
cos[9921]=78;
cos[9922]=78;
cos[9923]=78;
cos[9924]=78;
cos[9925]=78;
cos[9926]=78;
cos[9927]=78;
cos[9928]=78;
cos[9929]=78;
cos[9930]=78;
cos[9931]=78;
cos[9932]=78;
cos[9933]=78;
cos[9934]=78;
cos[9935]=78;
cos[9936]=78;
cos[9937]=78;
cos[9938]=78;
cos[9939]=78;
cos[9940]=78;
cos[9941]=78;
cos[9942]=78;
cos[9943]=78;
cos[9944]=78;
cos[9945]=78;
cos[9946]=78;
cos[9947]=78;
cos[9948]=78;
cos[9949]=78;
cos[9950]=78;
cos[9951]=78;
cos[9952]=78;
cos[9953]=78;
cos[9954]=78;
cos[9955]=78;
cos[9956]=78;
cos[9957]=78;
cos[9958]=78;
cos[9959]=78;
cos[9960]=78;
cos[9961]=78;
cos[9962]=78;
cos[9963]=78;
cos[9964]=78;
cos[9965]=78;
cos[9966]=78;
cos[9967]=78;
cos[9968]=78;
cos[9969]=78;
cos[9970]=78;
cos[9971]=78;
cos[9972]=78;
cos[9973]=78;
cos[9974]=78;
cos[9975]=78;
cos[9976]=78;
cos[9977]=78;
cos[9978]=78;
cos[9979]=78;
cos[9980]=78;
cos[9981]=78;
cos[9982]=78;
cos[9983]=78;
cos[9984]=78;
cos[9985]=78;
cos[9986]=78;
cos[9987]=78;
cos[9988]=78;
cos[9989]=78;
cos[9990]=78;
cos[9991]=78;
cos[9992]=78;
cos[9993]=78;
cos[9994]=78;
cos[9995]=78;
cos[9996]=78;
cos[9997]=78;
cos[9998]=78;
cos[9999]=78;
cos[10000]=78;
cos[10001]=78;
cos[10002]=78;
cos[10003]=78;
cos[10004]=78;
cos[10005]=78;
cos[10006]=78;
cos[10007]=78;
cos[10008]=78;
cos[10009]=78;
cos[10010]=78;
cos[10011]=78;
cos[10012]=78;
cos[10013]=78;
cos[10014]=78;
cos[10015]=78;
cos[10016]=78;
cos[10017]=78;
cos[10018]=78;
cos[10019]=78;
cos[10020]=78;
cos[10021]=78;
cos[10022]=78;
cos[10023]=78;
cos[10024]=78;
cos[10025]=78;
cos[10026]=78;
cos[10027]=78;
cos[10028]=78;
cos[10029]=78;
cos[10030]=78;
cos[10031]=78;
cos[10032]=78;
cos[10033]=78;
cos[10034]=78;
cos[10035]=78;
cos[10036]=78;
cos[10037]=78;
cos[10038]=78;
cos[10039]=78;
cos[10040]=78;
cos[10041]=78;
cos[10042]=78;
cos[10043]=78;
cos[10044]=78;
cos[10045]=78;
cos[10046]=78;
cos[10047]=78;
cos[10048]=78;
cos[10049]=78;
cos[10050]=78;
cos[10051]=78;
cos[10052]=78;
cos[10053]=78;
cos[10054]=78;
cos[10055]=78;
cos[10056]=78;
cos[10057]=78;
cos[10058]=78;
cos[10059]=78;
cos[10060]=78;
cos[10061]=78;
cos[10062]=78;
cos[10063]=78;
cos[10064]=78;
cos[10065]=78;
cos[10066]=78;
cos[10067]=78;
cos[10068]=78;
cos[10069]=78;
cos[10070]=78;
cos[10071]=78;
cos[10072]=78;
cos[10073]=78;
cos[10074]=78;
cos[10075]=78;
cos[10076]=78;
cos[10077]=78;
cos[10078]=78;
cos[10079]=78;
cos[10080]=78;
cos[10081]=78;
cos[10082]=78;
cos[10083]=78;
cos[10084]=78;
cos[10085]=78;
cos[10086]=78;
cos[10087]=78;
cos[10088]=78;
cos[10089]=78;
cos[10090]=78;
cos[10091]=78;
cos[10092]=78;
cos[10093]=78;
cos[10094]=78;
cos[10095]=78;
cos[10096]=78;
cos[10097]=78;
cos[10098]=78;
cos[10099]=78;
cos[10100]=78;
cos[10101]=78;
cos[10102]=78;
cos[10103]=78;
cos[10104]=78;
cos[10105]=78;
cos[10106]=78;
cos[10107]=78;
cos[10108]=78;
cos[10109]=78;
cos[10110]=78;
cos[10111]=78;
cos[10112]=78;
cos[10113]=78;
cos[10114]=78;
cos[10115]=78;
cos[10116]=78;
cos[10117]=78;
cos[10118]=78;
cos[10119]=78;
cos[10120]=78;
cos[10121]=78;
cos[10122]=78;
cos[10123]=78;
cos[10124]=78;
cos[10125]=78;
cos[10126]=78;
cos[10127]=78;
cos[10128]=78;
cos[10129]=78;
cos[10130]=78;
cos[10131]=78;
cos[10132]=78;
cos[10133]=78;
cos[10134]=78;
cos[10135]=78;
cos[10136]=78;
cos[10137]=78;
cos[10138]=78;
cos[10139]=78;
cos[10140]=78;
cos[10141]=78;
cos[10142]=78;
cos[10143]=78;
cos[10144]=78;
cos[10145]=78;
cos[10146]=78;
cos[10147]=78;
cos[10148]=78;
cos[10149]=78;
cos[10150]=78;
cos[10151]=78;
cos[10152]=78;
cos[10153]=78;
cos[10154]=78;
cos[10155]=78;
cos[10156]=78;
cos[10157]=78;
cos[10158]=78;
cos[10159]=78;
cos[10160]=78;
cos[10161]=78;
cos[10162]=78;
cos[10163]=78;
cos[10164]=78;
cos[10165]=78;
cos[10166]=78;
cos[10167]=78;
cos[10168]=78;
cos[10169]=78;
cos[10170]=78;
cos[10171]=78;
cos[10172]=78;
cos[10173]=78;
cos[10174]=78;
cos[10175]=78;
cos[10176]=78;
cos[10177]=78;
cos[10178]=78;
cos[10179]=78;
cos[10180]=78;
cos[10181]=78;
cos[10182]=78;
cos[10183]=78;
cos[10184]=78;
cos[10185]=78;
cos[10186]=78;
cos[10187]=78;
cos[10188]=78;
cos[10189]=78;
cos[10190]=78;
cos[10191]=78;
cos[10192]=78;
cos[10193]=78;
cos[10194]=78;
cos[10195]=78;
cos[10196]=78;
cos[10197]=78;
cos[10198]=78;
cos[10199]=78;
cos[10200]=78;
cos[10201]=78;
cos[10202]=77;
cos[10203]=77;
cos[10204]=77;
cos[10205]=77;
cos[10206]=77;
cos[10207]=77;
cos[10208]=77;
cos[10209]=77;
cos[10210]=77;
cos[10211]=77;
cos[10212]=77;
cos[10213]=77;
cos[10214]=77;
cos[10215]=77;
cos[10216]=77;
cos[10217]=77;
cos[10218]=77;
cos[10219]=77;
cos[10220]=77;
cos[10221]=77;
cos[10222]=77;
cos[10223]=77;
cos[10224]=77;
cos[10225]=77;
cos[10226]=77;
cos[10227]=77;
cos[10228]=77;
cos[10229]=77;
cos[10230]=77;
cos[10231]=77;
cos[10232]=77;
cos[10233]=77;
cos[10234]=77;
cos[10235]=77;
cos[10236]=77;
cos[10237]=77;
cos[10238]=77;
cos[10239]=77;
cos[10240]=77;
cos[10241]=77;
cos[10242]=77;
cos[10243]=77;
cos[10244]=77;
cos[10245]=77;
cos[10246]=77;
cos[10247]=77;
cos[10248]=77;
cos[10249]=77;
cos[10250]=77;
cos[10251]=77;
cos[10252]=77;
cos[10253]=77;
cos[10254]=77;
cos[10255]=77;
cos[10256]=77;
cos[10257]=77;
cos[10258]=77;
cos[10259]=77;
cos[10260]=77;
cos[10261]=77;
cos[10262]=77;
cos[10263]=77;
cos[10264]=77;
cos[10265]=77;
cos[10266]=77;
cos[10267]=77;
cos[10268]=77;
cos[10269]=77;
cos[10270]=77;
cos[10271]=77;
cos[10272]=77;
cos[10273]=77;
cos[10274]=77;
cos[10275]=77;
cos[10276]=77;
cos[10277]=77;
cos[10278]=77;
cos[10279]=77;
cos[10280]=77;
cos[10281]=77;
cos[10282]=77;
cos[10283]=77;
cos[10284]=77;
cos[10285]=77;
cos[10286]=77;
cos[10287]=77;
cos[10288]=77;
cos[10289]=77;
cos[10290]=77;
cos[10291]=77;
cos[10292]=77;
cos[10293]=77;
cos[10294]=77;
cos[10295]=77;
cos[10296]=77;
cos[10297]=77;
cos[10298]=77;
cos[10299]=77;
cos[10300]=77;
cos[10301]=77;
cos[10302]=77;
cos[10303]=77;
cos[10304]=77;
cos[10305]=77;
cos[10306]=77;
cos[10307]=77;
cos[10308]=77;
cos[10309]=77;
cos[10310]=77;
cos[10311]=77;
cos[10312]=77;
cos[10313]=77;
cos[10314]=77;
cos[10315]=77;
cos[10316]=77;
cos[10317]=77;
cos[10318]=77;
cos[10319]=77;
cos[10320]=77;
cos[10321]=77;
cos[10322]=77;
cos[10323]=77;
cos[10324]=77;
cos[10325]=77;
cos[10326]=76;
cos[10327]=76;
cos[10328]=76;
cos[10329]=76;
cos[10330]=76;
cos[10331]=76;
cos[10332]=76;
cos[10333]=76;
cos[10334]=76;
cos[10335]=76;
cos[10336]=76;
cos[10337]=76;
cos[10338]=76;
cos[10339]=76;
cos[10340]=76;
cos[10341]=76;
cos[10342]=76;
cos[10343]=76;
cos[10344]=76;
cos[10345]=76;
cos[10346]=76;
cos[10347]=76;
cos[10348]=76;
cos[10349]=76;
cos[10350]=76;
cos[10351]=76;
cos[10352]=76;
cos[10353]=76;
cos[10354]=76;
cos[10355]=76;
cos[10356]=76;
cos[10357]=76;
cos[10358]=76;
cos[10359]=76;
cos[10360]=76;
cos[10361]=76;
cos[10362]=76;
cos[10363]=76;
cos[10364]=76;
cos[10365]=76;
cos[10366]=76;
cos[10367]=76;
cos[10368]=76;
cos[10369]=76;
cos[10370]=76;
cos[10371]=76;
cos[10372]=76;
cos[10373]=76;
cos[10374]=76;
cos[10375]=76;
cos[10376]=76;
cos[10377]=76;
cos[10378]=76;
cos[10379]=76;
cos[10380]=76;
cos[10381]=76;
cos[10382]=76;
cos[10383]=76;
cos[10384]=76;
cos[10385]=76;
cos[10386]=76;
cos[10387]=76;
cos[10388]=76;
cos[10389]=76;
cos[10390]=76;
cos[10391]=76;
cos[10392]=76;
cos[10393]=76;
cos[10394]=76;
cos[10395]=76;
cos[10396]=76;
cos[10397]=76;
cos[10398]=76;
cos[10399]=76;
cos[10400]=76;
cos[10401]=76;
cos[10402]=76;
cos[10403]=76;
cos[10404]=76;
cos[10405]=76;
cos[10406]=76;
cos[10407]=76;
cos[10408]=76;
cos[10409]=76;
cos[10410]=76;
cos[10411]=76;
cos[10412]=76;
cos[10413]=76;
cos[10414]=75;
cos[10415]=75;
cos[10416]=75;
cos[10417]=75;
cos[10418]=75;
cos[10419]=75;
cos[10420]=75;
cos[10421]=75;
cos[10422]=75;
cos[10423]=75;
cos[10424]=75;
cos[10425]=75;
cos[10426]=75;
cos[10427]=75;
cos[10428]=75;
cos[10429]=75;
cos[10430]=75;
cos[10431]=75;
cos[10432]=75;
cos[10433]=75;
cos[10434]=75;
cos[10435]=75;
cos[10436]=75;
cos[10437]=75;
cos[10438]=75;
cos[10439]=75;
cos[10440]=75;
cos[10441]=75;
cos[10442]=75;
cos[10443]=75;
cos[10444]=75;
cos[10445]=75;
cos[10446]=75;
cos[10447]=75;
cos[10448]=75;
cos[10449]=75;
cos[10450]=75;
cos[10451]=75;
cos[10452]=75;
cos[10453]=75;
cos[10454]=75;
cos[10455]=75;
cos[10456]=75;
cos[10457]=75;
cos[10458]=75;
cos[10459]=75;
cos[10460]=75;
cos[10461]=75;
cos[10462]=75;
cos[10463]=75;
cos[10464]=75;
cos[10465]=75;
cos[10466]=75;
cos[10467]=75;
cos[10468]=75;
cos[10469]=75;
cos[10470]=75;
cos[10471]=75;
cos[10472]=75;
cos[10473]=75;
cos[10474]=75;
cos[10475]=75;
cos[10476]=75;
cos[10477]=75;
cos[10478]=75;
cos[10479]=75;
cos[10480]=75;
cos[10481]=75;
cos[10482]=75;
cos[10483]=75;
cos[10484]=75;
cos[10485]=75;
cos[10486]=75;
cos[10487]=74;
cos[10488]=74;
cos[10489]=74;
cos[10490]=74;
cos[10491]=74;
cos[10492]=74;
cos[10493]=74;
cos[10494]=74;
cos[10495]=74;
cos[10496]=74;
cos[10497]=74;
cos[10498]=74;
cos[10499]=74;
cos[10500]=74;
cos[10501]=74;
cos[10502]=74;
cos[10503]=74;
cos[10504]=74;
cos[10505]=74;
cos[10506]=74;
cos[10507]=74;
cos[10508]=74;
cos[10509]=74;
cos[10510]=74;
cos[10511]=74;
cos[10512]=74;
cos[10513]=74;
cos[10514]=74;
cos[10515]=74;
cos[10516]=74;
cos[10517]=74;
cos[10518]=74;
cos[10519]=74;
cos[10520]=74;
cos[10521]=74;
cos[10522]=74;
cos[10523]=74;
cos[10524]=74;
cos[10525]=74;
cos[10526]=74;
cos[10527]=74;
cos[10528]=74;
cos[10529]=74;
cos[10530]=74;
cos[10531]=74;
cos[10532]=74;
cos[10533]=74;
cos[10534]=74;
cos[10535]=74;
cos[10536]=74;
cos[10537]=74;
cos[10538]=74;
cos[10539]=74;
cos[10540]=74;
cos[10541]=74;
cos[10542]=74;
cos[10543]=74;
cos[10544]=74;
cos[10545]=74;
cos[10546]=74;
cos[10547]=74;
cos[10548]=74;
cos[10549]=74;
cos[10550]=74;
cos[10551]=73;
cos[10552]=73;
cos[10553]=73;
cos[10554]=73;
cos[10555]=73;
cos[10556]=73;
cos[10557]=73;
cos[10558]=73;
cos[10559]=73;
cos[10560]=73;
cos[10561]=73;
cos[10562]=73;
cos[10563]=73;
cos[10564]=73;
cos[10565]=73;
cos[10566]=73;
cos[10567]=73;
cos[10568]=73;
cos[10569]=73;
cos[10570]=73;
cos[10571]=73;
cos[10572]=73;
cos[10573]=73;
cos[10574]=73;
cos[10575]=73;
cos[10576]=73;
cos[10577]=73;
cos[10578]=73;
cos[10579]=73;
cos[10580]=73;
cos[10581]=73;
cos[10582]=73;
cos[10583]=73;
cos[10584]=73;
cos[10585]=73;
cos[10586]=73;
cos[10587]=73;
cos[10588]=73;
cos[10589]=73;
cos[10590]=73;
cos[10591]=73;
cos[10592]=73;
cos[10593]=73;
cos[10594]=73;
cos[10595]=73;
cos[10596]=73;
cos[10597]=73;
cos[10598]=73;
cos[10599]=73;
cos[10600]=73;
cos[10601]=73;
cos[10602]=73;
cos[10603]=73;
cos[10604]=73;
cos[10605]=73;
cos[10606]=73;
cos[10607]=73;
cos[10608]=72;
cos[10609]=72;
cos[10610]=72;
cos[10611]=72;
cos[10612]=72;
cos[10613]=72;
cos[10614]=72;
cos[10615]=72;
cos[10616]=72;
cos[10617]=72;
cos[10618]=72;
cos[10619]=72;
cos[10620]=72;
cos[10621]=72;
cos[10622]=72;
cos[10623]=72;
cos[10624]=72;
cos[10625]=72;
cos[10626]=72;
cos[10627]=72;
cos[10628]=72;
cos[10629]=72;
cos[10630]=72;
cos[10631]=72;
cos[10632]=72;
cos[10633]=72;
cos[10634]=72;
cos[10635]=72;
cos[10636]=72;
cos[10637]=72;
cos[10638]=72;
cos[10639]=72;
cos[10640]=72;
cos[10641]=72;
cos[10642]=72;
cos[10643]=72;
cos[10644]=72;
cos[10645]=72;
cos[10646]=72;
cos[10647]=72;
cos[10648]=72;
cos[10649]=72;
cos[10650]=72;
cos[10651]=72;
cos[10652]=72;
cos[10653]=72;
cos[10654]=72;
cos[10655]=72;
cos[10656]=72;
cos[10657]=72;
cos[10658]=72;
cos[10659]=72;
cos[10660]=72;
cos[10661]=71;
cos[10662]=71;
cos[10663]=71;
cos[10664]=71;
cos[10665]=71;
cos[10666]=71;
cos[10667]=71;
cos[10668]=71;
cos[10669]=71;
cos[10670]=71;
cos[10671]=71;
cos[10672]=71;
cos[10673]=71;
cos[10674]=71;
cos[10675]=71;
cos[10676]=71;
cos[10677]=71;
cos[10678]=71;
cos[10679]=71;
cos[10680]=71;
cos[10681]=71;
cos[10682]=71;
cos[10683]=71;
cos[10684]=71;
cos[10685]=71;
cos[10686]=71;
cos[10687]=71;
cos[10688]=71;
cos[10689]=71;
cos[10690]=71;
cos[10691]=71;
cos[10692]=71;
cos[10693]=71;
cos[10694]=71;
cos[10695]=71;
cos[10696]=71;
cos[10697]=71;
cos[10698]=71;
cos[10699]=71;
cos[10700]=71;
cos[10701]=71;
cos[10702]=71;
cos[10703]=71;
cos[10704]=71;
cos[10705]=71;
cos[10706]=71;
cos[10707]=71;
cos[10708]=71;
cos[10709]=71;
cos[10710]=70;
cos[10711]=70;
cos[10712]=70;
cos[10713]=70;
cos[10714]=70;
cos[10715]=70;
cos[10716]=70;
cos[10717]=70;
cos[10718]=70;
cos[10719]=70;
cos[10720]=70;
cos[10721]=70;
cos[10722]=70;
cos[10723]=70;
cos[10724]=70;
cos[10725]=70;
cos[10726]=70;
cos[10727]=70;
cos[10728]=70;
cos[10729]=70;
cos[10730]=70;
cos[10731]=70;
cos[10732]=70;
cos[10733]=70;
cos[10734]=70;
cos[10735]=70;
cos[10736]=70;
cos[10737]=70;
cos[10738]=70;
cos[10739]=70;
cos[10740]=70;
cos[10741]=70;
cos[10742]=70;
cos[10743]=70;
cos[10744]=70;
cos[10745]=70;
cos[10746]=70;
cos[10747]=70;
cos[10748]=70;
cos[10749]=70;
cos[10750]=70;
cos[10751]=70;
cos[10752]=70;
cos[10753]=70;
cos[10754]=70;
cos[10755]=69;
cos[10756]=69;
cos[10757]=69;
cos[10758]=69;
cos[10759]=69;
cos[10760]=69;
cos[10761]=69;
cos[10762]=69;
cos[10763]=69;
cos[10764]=69;
cos[10765]=69;
cos[10766]=69;
cos[10767]=69;
cos[10768]=69;
cos[10769]=69;
cos[10770]=69;
cos[10771]=69;
cos[10772]=69;
cos[10773]=69;
cos[10774]=69;
cos[10775]=69;
cos[10776]=69;
cos[10777]=69;
cos[10778]=69;
cos[10779]=69;
cos[10780]=69;
cos[10781]=69;
cos[10782]=69;
cos[10783]=69;
cos[10784]=69;
cos[10785]=69;
cos[10786]=69;
cos[10787]=69;
cos[10788]=69;
cos[10789]=69;
cos[10790]=69;
cos[10791]=69;
cos[10792]=69;
cos[10793]=69;
cos[10794]=69;
cos[10795]=69;
cos[10796]=69;
cos[10797]=69;
cos[10798]=69;
cos[10799]=68;
cos[10800]=68;
cos[10801]=68;
cos[10802]=68;
cos[10803]=68;
cos[10804]=68;
cos[10805]=68;
cos[10806]=68;
cos[10807]=68;
cos[10808]=68;
cos[10809]=68;
cos[10810]=68;
cos[10811]=68;
cos[10812]=68;
cos[10813]=68;
cos[10814]=68;
cos[10815]=68;
cos[10816]=68;
cos[10817]=68;
cos[10818]=68;
cos[10819]=68;
cos[10820]=68;
cos[10821]=68;
cos[10822]=68;
cos[10823]=68;
cos[10824]=68;
cos[10825]=68;
cos[10826]=68;
cos[10827]=68;
cos[10828]=68;
cos[10829]=68;
cos[10830]=68;
cos[10831]=68;
cos[10832]=68;
cos[10833]=68;
cos[10834]=68;
cos[10835]=68;
cos[10836]=68;
cos[10837]=68;
cos[10838]=68;
cos[10839]=68;
cos[10840]=67;
cos[10841]=67;
cos[10842]=67;
cos[10843]=67;
cos[10844]=67;
cos[10845]=67;
cos[10846]=67;
cos[10847]=67;
cos[10848]=67;
cos[10849]=67;
cos[10850]=67;
cos[10851]=67;
cos[10852]=67;
cos[10853]=67;
cos[10854]=67;
cos[10855]=67;
cos[10856]=67;
cos[10857]=67;
cos[10858]=67;
cos[10859]=67;
cos[10860]=67;
cos[10861]=67;
cos[10862]=67;
cos[10863]=67;
cos[10864]=67;
cos[10865]=67;
cos[10866]=67;
cos[10867]=67;
cos[10868]=67;
cos[10869]=67;
cos[10870]=67;
cos[10871]=67;
cos[10872]=67;
cos[10873]=67;
cos[10874]=67;
cos[10875]=67;
cos[10876]=67;
cos[10877]=67;
cos[10878]=67;
cos[10879]=67;
cos[10880]=66;
cos[10881]=66;
cos[10882]=66;
cos[10883]=66;
cos[10884]=66;
cos[10885]=66;
cos[10886]=66;
cos[10887]=66;
cos[10888]=66;
cos[10889]=66;
cos[10890]=66;
cos[10891]=66;
cos[10892]=66;
cos[10893]=66;
cos[10894]=66;
cos[10895]=66;
cos[10896]=66;
cos[10897]=66;
cos[10898]=66;
cos[10899]=66;
cos[10900]=66;
cos[10901]=66;
cos[10902]=66;
cos[10903]=66;
cos[10904]=66;
cos[10905]=66;
cos[10906]=66;
cos[10907]=66;
cos[10908]=66;
cos[10909]=66;
cos[10910]=66;
cos[10911]=66;
cos[10912]=66;
cos[10913]=66;
cos[10914]=66;
cos[10915]=66;
cos[10916]=66;
cos[10917]=66;
cos[10918]=65;
cos[10919]=65;
cos[10920]=65;
cos[10921]=65;
cos[10922]=65;
cos[10923]=65;
cos[10924]=65;
cos[10925]=65;
cos[10926]=65;
cos[10927]=65;
cos[10928]=65;
cos[10929]=65;
cos[10930]=65;
cos[10931]=65;
cos[10932]=65;
cos[10933]=65;
cos[10934]=65;
cos[10935]=65;
cos[10936]=65;
cos[10937]=65;
cos[10938]=65;
cos[10939]=65;
cos[10940]=65;
cos[10941]=65;
cos[10942]=65;
cos[10943]=65;
cos[10944]=65;
cos[10945]=65;
cos[10946]=65;
cos[10947]=65;
cos[10948]=65;
cos[10949]=65;
cos[10950]=65;
cos[10951]=65;
cos[10952]=65;
cos[10953]=65;
cos[10954]=65;
cos[10955]=64;
cos[10956]=64;
cos[10957]=64;
cos[10958]=64;
cos[10959]=64;
cos[10960]=64;
cos[10961]=64;
cos[10962]=64;
cos[10963]=64;
cos[10964]=64;
cos[10965]=64;
cos[10966]=64;
cos[10967]=64;
cos[10968]=64;
cos[10969]=64;
cos[10970]=64;
cos[10971]=64;
cos[10972]=64;
cos[10973]=64;
cos[10974]=64;
cos[10975]=64;
cos[10976]=64;
cos[10977]=64;
cos[10978]=64;
cos[10979]=64;
cos[10980]=64;
cos[10981]=64;
cos[10982]=64;
cos[10983]=64;
cos[10984]=64;
cos[10985]=64;
cos[10986]=64;
cos[10987]=64;
cos[10988]=64;
cos[10989]=64;
cos[10990]=63;
cos[10991]=63;
cos[10992]=63;
cos[10993]=63;
cos[10994]=63;
cos[10995]=63;
cos[10996]=63;
cos[10997]=63;
cos[10998]=63;
cos[10999]=63;
cos[11000]=63;
cos[11001]=63;
cos[11002]=63;
cos[11003]=63;
cos[11004]=63;
cos[11005]=63;
cos[11006]=63;
cos[11007]=63;
cos[11008]=63;
cos[11009]=63;
cos[11010]=63;
cos[11011]=63;
cos[11012]=63;
cos[11013]=63;
cos[11014]=63;
cos[11015]=63;
cos[11016]=63;
cos[11017]=63;
cos[11018]=63;
cos[11019]=63;
cos[11020]=63;
cos[11021]=63;
cos[11022]=63;
cos[11023]=63;
cos[11024]=63;
cos[11025]=62;
cos[11026]=62;
cos[11027]=62;
cos[11028]=62;
cos[11029]=62;
cos[11030]=62;
cos[11031]=62;
cos[11032]=62;
cos[11033]=62;
cos[11034]=62;
cos[11035]=62;
cos[11036]=62;
cos[11037]=62;
cos[11038]=62;
cos[11039]=62;
cos[11040]=62;
cos[11041]=62;
cos[11042]=62;
cos[11043]=62;
cos[11044]=62;
cos[11045]=62;
cos[11046]=62;
cos[11047]=62;
cos[11048]=62;
cos[11049]=62;
cos[11050]=62;
cos[11051]=62;
cos[11052]=62;
cos[11053]=62;
cos[11054]=62;
cos[11055]=62;
cos[11056]=62;
cos[11057]=62;
cos[11058]=61;
cos[11059]=61;
cos[11060]=61;
cos[11061]=61;
cos[11062]=61;
cos[11063]=61;
cos[11064]=61;
cos[11065]=61;
cos[11066]=61;
cos[11067]=61;
cos[11068]=61;
cos[11069]=61;
cos[11070]=61;
cos[11071]=61;
cos[11072]=61;
cos[11073]=61;
cos[11074]=61;
cos[11075]=61;
cos[11076]=61;
cos[11077]=61;
cos[11078]=61;
cos[11079]=61;
cos[11080]=61;
cos[11081]=61;
cos[11082]=61;
cos[11083]=61;
cos[11084]=61;
cos[11085]=61;
cos[11086]=61;
cos[11087]=61;
cos[11088]=61;
cos[11089]=61;
cos[11090]=61;
cos[11091]=60;
cos[11092]=60;
cos[11093]=60;
cos[11094]=60;
cos[11095]=60;
cos[11096]=60;
cos[11097]=60;
cos[11098]=60;
cos[11099]=60;
cos[11100]=60;
cos[11101]=60;
cos[11102]=60;
cos[11103]=60;
cos[11104]=60;
cos[11105]=60;
cos[11106]=60;
cos[11107]=60;
cos[11108]=60;
cos[11109]=60;
cos[11110]=60;
cos[11111]=60;
cos[11112]=60;
cos[11113]=60;
cos[11114]=60;
cos[11115]=60;
cos[11116]=60;
cos[11117]=60;
cos[11118]=60;
cos[11119]=60;
cos[11120]=60;
cos[11121]=60;
cos[11122]=60;
cos[11123]=59;
cos[11124]=59;
cos[11125]=59;
cos[11126]=59;
cos[11127]=59;
cos[11128]=59;
cos[11129]=59;
cos[11130]=59;
cos[11131]=59;
cos[11132]=59;
cos[11133]=59;
cos[11134]=59;
cos[11135]=59;
cos[11136]=59;
cos[11137]=59;
cos[11138]=59;
cos[11139]=59;
cos[11140]=59;
cos[11141]=59;
cos[11142]=59;
cos[11143]=59;
cos[11144]=59;
cos[11145]=59;
cos[11146]=59;
cos[11147]=59;
cos[11148]=59;
cos[11149]=59;
cos[11150]=59;
cos[11151]=59;
cos[11152]=59;
cos[11153]=59;
cos[11154]=58;
cos[11155]=58;
cos[11156]=58;
cos[11157]=58;
cos[11158]=58;
cos[11159]=58;
cos[11160]=58;
cos[11161]=58;
cos[11162]=58;
cos[11163]=58;
cos[11164]=58;
cos[11165]=58;
cos[11166]=58;
cos[11167]=58;
cos[11168]=58;
cos[11169]=58;
cos[11170]=58;
cos[11171]=58;
cos[11172]=58;
cos[11173]=58;
cos[11174]=58;
cos[11175]=58;
cos[11176]=58;
cos[11177]=58;
cos[11178]=58;
cos[11179]=58;
cos[11180]=58;
cos[11181]=58;
cos[11182]=58;
cos[11183]=58;
cos[11184]=57;
cos[11185]=57;
cos[11186]=57;
cos[11187]=57;
cos[11188]=57;
cos[11189]=57;
cos[11190]=57;
cos[11191]=57;
cos[11192]=57;
cos[11193]=57;
cos[11194]=57;
cos[11195]=57;
cos[11196]=57;
cos[11197]=57;
cos[11198]=57;
cos[11199]=57;
cos[11200]=57;
cos[11201]=57;
cos[11202]=57;
cos[11203]=57;
cos[11204]=57;
cos[11205]=57;
cos[11206]=57;
cos[11207]=57;
cos[11208]=57;
cos[11209]=57;
cos[11210]=57;
cos[11211]=57;
cos[11212]=57;
cos[11213]=57;
cos[11214]=56;
cos[11215]=56;
cos[11216]=56;
cos[11217]=56;
cos[11218]=56;
cos[11219]=56;
cos[11220]=56;
cos[11221]=56;
cos[11222]=56;
cos[11223]=56;
cos[11224]=56;
cos[11225]=56;
cos[11226]=56;
cos[11227]=56;
cos[11228]=56;
cos[11229]=56;
cos[11230]=56;
cos[11231]=56;
cos[11232]=56;
cos[11233]=56;
cos[11234]=56;
cos[11235]=56;
cos[11236]=56;
cos[11237]=56;
cos[11238]=56;
cos[11239]=56;
cos[11240]=56;
cos[11241]=56;
cos[11242]=56;
cos[11243]=55;
cos[11244]=55;
cos[11245]=55;
cos[11246]=55;
cos[11247]=55;
cos[11248]=55;
cos[11249]=55;
cos[11250]=55;
cos[11251]=55;
cos[11252]=55;
cos[11253]=55;
cos[11254]=55;
cos[11255]=55;
cos[11256]=55;
cos[11257]=55;
cos[11258]=55;
cos[11259]=55;
cos[11260]=55;
cos[11261]=55;
cos[11262]=55;
cos[11263]=55;
cos[11264]=55;
cos[11265]=55;
cos[11266]=55;
cos[11267]=55;
cos[11268]=55;
cos[11269]=55;
cos[11270]=55;
cos[11271]=55;
cos[11272]=54;
cos[11273]=54;
cos[11274]=54;
cos[11275]=54;
cos[11276]=54;
cos[11277]=54;
cos[11278]=54;
cos[11279]=54;
cos[11280]=54;
cos[11281]=54;
cos[11282]=54;
cos[11283]=54;
cos[11284]=54;
cos[11285]=54;
cos[11286]=54;
cos[11287]=54;
cos[11288]=54;
cos[11289]=54;
cos[11290]=54;
cos[11291]=54;
cos[11292]=54;
cos[11293]=54;
cos[11294]=54;
cos[11295]=54;
cos[11296]=54;
cos[11297]=54;
cos[11298]=54;
cos[11299]=54;
cos[11300]=53;
cos[11301]=53;
cos[11302]=53;
cos[11303]=53;
cos[11304]=53;
cos[11305]=53;
cos[11306]=53;
cos[11307]=53;
cos[11308]=53;
cos[11309]=53;
cos[11310]=53;
cos[11311]=53;
cos[11312]=53;
cos[11313]=53;
cos[11314]=53;
cos[11315]=53;
cos[11316]=53;
cos[11317]=53;
cos[11318]=53;
cos[11319]=53;
cos[11320]=53;
cos[11321]=53;
cos[11322]=53;
cos[11323]=53;
cos[11324]=53;
cos[11325]=53;
cos[11326]=53;
cos[11327]=53;
cos[11328]=52;
cos[11329]=52;
cos[11330]=52;
cos[11331]=52;
cos[11332]=52;
cos[11333]=52;
cos[11334]=52;
cos[11335]=52;
cos[11336]=52;
cos[11337]=52;
cos[11338]=52;
cos[11339]=52;
cos[11340]=52;
cos[11341]=52;
cos[11342]=52;
cos[11343]=52;
cos[11344]=52;
cos[11345]=52;
cos[11346]=52;
cos[11347]=52;
cos[11348]=52;
cos[11349]=52;
cos[11350]=52;
cos[11351]=52;
cos[11352]=52;
cos[11353]=52;
cos[11354]=52;
cos[11355]=51;
cos[11356]=51;
cos[11357]=51;
cos[11358]=51;
cos[11359]=51;
cos[11360]=51;
cos[11361]=51;
cos[11362]=51;
cos[11363]=51;
cos[11364]=51;
cos[11365]=51;
cos[11366]=51;
cos[11367]=51;
cos[11368]=51;
cos[11369]=51;
cos[11370]=51;
cos[11371]=51;
cos[11372]=51;
cos[11373]=51;
cos[11374]=51;
cos[11375]=51;
cos[11376]=51;
cos[11377]=51;
cos[11378]=51;
cos[11379]=51;
cos[11380]=51;
cos[11381]=51;
cos[11382]=50;
cos[11383]=50;
cos[11384]=50;
cos[11385]=50;
cos[11386]=50;
cos[11387]=50;
cos[11388]=50;
cos[11389]=50;
cos[11390]=50;
cos[11391]=50;
cos[11392]=50;
cos[11393]=50;
cos[11394]=50;
cos[11395]=50;
cos[11396]=50;
cos[11397]=50;
cos[11398]=50;
cos[11399]=50;
cos[11400]=50;
cos[11401]=50;
cos[11402]=50;
cos[11403]=50;
cos[11404]=50;
cos[11405]=50;
cos[11406]=50;
cos[11407]=50;
cos[11408]=49;
cos[11409]=49;
cos[11410]=49;
cos[11411]=49;
cos[11412]=49;
cos[11413]=49;
cos[11414]=49;
cos[11415]=49;
cos[11416]=49;
cos[11417]=49;
cos[11418]=49;
cos[11419]=49;
cos[11420]=49;
cos[11421]=49;
cos[11422]=49;
cos[11423]=49;
cos[11424]=49;
cos[11425]=49;
cos[11426]=49;
cos[11427]=49;
cos[11428]=49;
cos[11429]=49;
cos[11430]=49;
cos[11431]=49;
cos[11432]=49;
cos[11433]=49;
cos[11434]=49;
cos[11435]=48;
cos[11436]=48;
cos[11437]=48;
cos[11438]=48;
cos[11439]=48;
cos[11440]=48;
cos[11441]=48;
cos[11442]=48;
cos[11443]=48;
cos[11444]=48;
cos[11445]=48;
cos[11446]=48;
cos[11447]=48;
cos[11448]=48;
cos[11449]=48;
cos[11450]=48;
cos[11451]=48;
cos[11452]=48;
cos[11453]=48;
cos[11454]=48;
cos[11455]=48;
cos[11456]=48;
cos[11457]=48;
cos[11458]=48;
cos[11459]=48;
cos[11460]=47;
cos[11461]=47;
cos[11462]=47;
cos[11463]=47;
cos[11464]=47;
cos[11465]=47;
cos[11466]=47;
cos[11467]=47;
cos[11468]=47;
cos[11469]=47;
cos[11470]=47;
cos[11471]=47;
cos[11472]=47;
cos[11473]=47;
cos[11474]=47;
cos[11475]=47;
cos[11476]=47;
cos[11477]=47;
cos[11478]=47;
cos[11479]=47;
cos[11480]=47;
cos[11481]=47;
cos[11482]=47;
cos[11483]=47;
cos[11484]=47;
cos[11485]=47;
cos[11486]=46;
cos[11487]=46;
cos[11488]=46;
cos[11489]=46;
cos[11490]=46;
cos[11491]=46;
cos[11492]=46;
cos[11493]=46;
cos[11494]=46;
cos[11495]=46;
cos[11496]=46;
cos[11497]=46;
cos[11498]=46;
cos[11499]=46;
cos[11500]=46;
cos[11501]=46;
cos[11502]=46;
cos[11503]=46;
cos[11504]=46;
cos[11505]=46;
cos[11506]=46;
cos[11507]=46;
cos[11508]=46;
cos[11509]=46;
cos[11510]=46;
cos[11511]=45;
cos[11512]=45;
cos[11513]=45;
cos[11514]=45;
cos[11515]=45;
cos[11516]=45;
cos[11517]=45;
cos[11518]=45;
cos[11519]=45;
cos[11520]=45;
cos[11521]=45;
cos[11522]=45;
cos[11523]=45;
cos[11524]=45;
cos[11525]=45;
cos[11526]=45;
cos[11527]=45;
cos[11528]=45;
cos[11529]=45;
cos[11530]=45;
cos[11531]=45;
cos[11532]=45;
cos[11533]=45;
cos[11534]=45;
cos[11535]=45;
cos[11536]=44;
cos[11537]=44;
cos[11538]=44;
cos[11539]=44;
cos[11540]=44;
cos[11541]=44;
cos[11542]=44;
cos[11543]=44;
cos[11544]=44;
cos[11545]=44;
cos[11546]=44;
cos[11547]=44;
cos[11548]=44;
cos[11549]=44;
cos[11550]=44;
cos[11551]=44;
cos[11552]=44;
cos[11553]=44;
cos[11554]=44;
cos[11555]=44;
cos[11556]=44;
cos[11557]=44;
cos[11558]=44;
cos[11559]=44;
cos[11560]=44;
cos[11561]=43;
cos[11562]=43;
cos[11563]=43;
cos[11564]=43;
cos[11565]=43;
cos[11566]=43;
cos[11567]=43;
cos[11568]=43;
cos[11569]=43;
cos[11570]=43;
cos[11571]=43;
cos[11572]=43;
cos[11573]=43;
cos[11574]=43;
cos[11575]=43;
cos[11576]=43;
cos[11577]=43;
cos[11578]=43;
cos[11579]=43;
cos[11580]=43;
cos[11581]=43;
cos[11582]=43;
cos[11583]=43;
cos[11584]=43;
cos[11585]=42;
cos[11586]=42;
cos[11587]=42;
cos[11588]=42;
cos[11589]=42;
cos[11590]=42;
cos[11591]=42;
cos[11592]=42;
cos[11593]=42;
cos[11594]=42;
cos[11595]=42;
cos[11596]=42;
cos[11597]=42;
cos[11598]=42;
cos[11599]=42;
cos[11600]=42;
cos[11601]=42;
cos[11602]=42;
cos[11603]=42;
cos[11604]=42;
cos[11605]=42;
cos[11606]=42;
cos[11607]=42;
cos[11608]=42;
cos[11609]=41;
cos[11610]=41;
cos[11611]=41;
cos[11612]=41;
cos[11613]=41;
cos[11614]=41;
cos[11615]=41;
cos[11616]=41;
cos[11617]=41;
cos[11618]=41;
cos[11619]=41;
cos[11620]=41;
cos[11621]=41;
cos[11622]=41;
cos[11623]=41;
cos[11624]=41;
cos[11625]=41;
cos[11626]=41;
cos[11627]=41;
cos[11628]=41;
cos[11629]=41;
cos[11630]=41;
cos[11631]=41;
cos[11632]=41;
cos[11633]=40;
cos[11634]=40;
cos[11635]=40;
cos[11636]=40;
cos[11637]=40;
cos[11638]=40;
cos[11639]=40;
cos[11640]=40;
cos[11641]=40;
cos[11642]=40;
cos[11643]=40;
cos[11644]=40;
cos[11645]=40;
cos[11646]=40;
cos[11647]=40;
cos[11648]=40;
cos[11649]=40;
cos[11650]=40;
cos[11651]=40;
cos[11652]=40;
cos[11653]=40;
cos[11654]=40;
cos[11655]=40;
cos[11656]=40;
cos[11657]=39;
cos[11658]=39;
cos[11659]=39;
cos[11660]=39;
cos[11661]=39;
cos[11662]=39;
cos[11663]=39;
cos[11664]=39;
cos[11665]=39;
cos[11666]=39;
cos[11667]=39;
cos[11668]=39;
cos[11669]=39;
cos[11670]=39;
cos[11671]=39;
cos[11672]=39;
cos[11673]=39;
cos[11674]=39;
cos[11675]=39;
cos[11676]=39;
cos[11677]=39;
cos[11678]=39;
cos[11679]=39;
cos[11680]=38;
cos[11681]=38;
cos[11682]=38;
cos[11683]=38;
cos[11684]=38;
cos[11685]=38;
cos[11686]=38;
cos[11687]=38;
cos[11688]=38;
cos[11689]=38;
cos[11690]=38;
cos[11691]=38;
cos[11692]=38;
cos[11693]=38;
cos[11694]=38;
cos[11695]=38;
cos[11696]=38;
cos[11697]=38;
cos[11698]=38;
cos[11699]=38;
cos[11700]=38;
cos[11701]=38;
cos[11702]=38;
cos[11703]=38;
cos[11704]=37;
cos[11705]=37;
cos[11706]=37;
cos[11707]=37;
cos[11708]=37;
cos[11709]=37;
cos[11710]=37;
cos[11711]=37;
cos[11712]=37;
cos[11713]=37;
cos[11714]=37;
cos[11715]=37;
cos[11716]=37;
cos[11717]=37;
cos[11718]=37;
cos[11719]=37;
cos[11720]=37;
cos[11721]=37;
cos[11722]=37;
cos[11723]=37;
cos[11724]=37;
cos[11725]=37;
cos[11726]=37;
cos[11727]=36;
cos[11728]=36;
cos[11729]=36;
cos[11730]=36;
cos[11731]=36;
cos[11732]=36;
cos[11733]=36;
cos[11734]=36;
cos[11735]=36;
cos[11736]=36;
cos[11737]=36;
cos[11738]=36;
cos[11739]=36;
cos[11740]=36;
cos[11741]=36;
cos[11742]=36;
cos[11743]=36;
cos[11744]=36;
cos[11745]=36;
cos[11746]=36;
cos[11747]=36;
cos[11748]=36;
cos[11749]=36;
cos[11750]=35;
cos[11751]=35;
cos[11752]=35;
cos[11753]=35;
cos[11754]=35;
cos[11755]=35;
cos[11756]=35;
cos[11757]=35;
cos[11758]=35;
cos[11759]=35;
cos[11760]=35;
cos[11761]=35;
cos[11762]=35;
cos[11763]=35;
cos[11764]=35;
cos[11765]=35;
cos[11766]=35;
cos[11767]=35;
cos[11768]=35;
cos[11769]=35;
cos[11770]=35;
cos[11771]=35;
cos[11772]=35;
cos[11773]=34;
cos[11774]=34;
cos[11775]=34;
cos[11776]=34;
cos[11777]=34;
cos[11778]=34;
cos[11779]=34;
cos[11780]=34;
cos[11781]=34;
cos[11782]=34;
cos[11783]=34;
cos[11784]=34;
cos[11785]=34;
cos[11786]=34;
cos[11787]=34;
cos[11788]=34;
cos[11789]=34;
cos[11790]=34;
cos[11791]=34;
cos[11792]=34;
cos[11793]=34;
cos[11794]=34;
cos[11795]=33;
cos[11796]=33;
cos[11797]=33;
cos[11798]=33;
cos[11799]=33;
cos[11800]=33;
cos[11801]=33;
cos[11802]=33;
cos[11803]=33;
cos[11804]=33;
cos[11805]=33;
cos[11806]=33;
cos[11807]=33;
cos[11808]=33;
cos[11809]=33;
cos[11810]=33;
cos[11811]=33;
cos[11812]=33;
cos[11813]=33;
cos[11814]=33;
cos[11815]=33;
cos[11816]=33;
cos[11817]=33;
cos[11818]=32;
cos[11819]=32;
cos[11820]=32;
cos[11821]=32;
cos[11822]=32;
cos[11823]=32;
cos[11824]=32;
cos[11825]=32;
cos[11826]=32;
cos[11827]=32;
cos[11828]=32;
cos[11829]=32;
cos[11830]=32;
cos[11831]=32;
cos[11832]=32;
cos[11833]=32;
cos[11834]=32;
cos[11835]=32;
cos[11836]=32;
cos[11837]=32;
cos[11838]=32;
cos[11839]=32;
cos[11840]=31;
cos[11841]=31;
cos[11842]=31;
cos[11843]=31;
cos[11844]=31;
cos[11845]=31;
cos[11846]=31;
cos[11847]=31;
cos[11848]=31;
cos[11849]=31;
cos[11850]=31;
cos[11851]=31;
cos[11852]=31;
cos[11853]=31;
cos[11854]=31;
cos[11855]=31;
cos[11856]=31;
cos[11857]=31;
cos[11858]=31;
cos[11859]=31;
cos[11860]=31;
cos[11861]=31;
cos[11862]=30;
cos[11863]=30;
cos[11864]=30;
cos[11865]=30;
cos[11866]=30;
cos[11867]=30;
cos[11868]=30;
cos[11869]=30;
cos[11870]=30;
cos[11871]=30;
cos[11872]=30;
cos[11873]=30;
cos[11874]=30;
cos[11875]=30;
cos[11876]=30;
cos[11877]=30;
cos[11878]=30;
cos[11879]=30;
cos[11880]=30;
cos[11881]=30;
cos[11882]=30;
cos[11883]=30;
cos[11884]=29;
cos[11885]=29;
cos[11886]=29;
cos[11887]=29;
cos[11888]=29;
cos[11889]=29;
cos[11890]=29;
cos[11891]=29;
cos[11892]=29;
cos[11893]=29;
cos[11894]=29;
cos[11895]=29;
cos[11896]=29;
cos[11897]=29;
cos[11898]=29;
cos[11899]=29;
cos[11900]=29;
cos[11901]=29;
cos[11902]=29;
cos[11903]=29;
cos[11904]=29;
cos[11905]=29;
cos[11906]=28;
cos[11907]=28;
cos[11908]=28;
cos[11909]=28;
cos[11910]=28;
cos[11911]=28;
cos[11912]=28;
cos[11913]=28;
cos[11914]=28;
cos[11915]=28;
cos[11916]=28;
cos[11917]=28;
cos[11918]=28;
cos[11919]=28;
cos[11920]=28;
cos[11921]=28;
cos[11922]=28;
cos[11923]=28;
cos[11924]=28;
cos[11925]=28;
cos[11926]=28;
cos[11927]=28;
cos[11928]=27;
cos[11929]=27;
cos[11930]=27;
cos[11931]=27;
cos[11932]=27;
cos[11933]=27;
cos[11934]=27;
cos[11935]=27;
cos[11936]=27;
cos[11937]=27;
cos[11938]=27;
cos[11939]=27;
cos[11940]=27;
cos[11941]=27;
cos[11942]=27;
cos[11943]=27;
cos[11944]=27;
cos[11945]=27;
cos[11946]=27;
cos[11947]=27;
cos[11948]=27;
cos[11949]=27;
cos[11950]=26;
cos[11951]=26;
cos[11952]=26;
cos[11953]=26;
cos[11954]=26;
cos[11955]=26;
cos[11956]=26;
cos[11957]=26;
cos[11958]=26;
cos[11959]=26;
cos[11960]=26;
cos[11961]=26;
cos[11962]=26;
cos[11963]=26;
cos[11964]=26;
cos[11965]=26;
cos[11966]=26;
cos[11967]=26;
cos[11968]=26;
cos[11969]=26;
cos[11970]=26;
cos[11971]=25;
cos[11972]=25;
cos[11973]=25;
cos[11974]=25;
cos[11975]=25;
cos[11976]=25;
cos[11977]=25;
cos[11978]=25;
cos[11979]=25;
cos[11980]=25;
cos[11981]=25;
cos[11982]=25;
cos[11983]=25;
cos[11984]=25;
cos[11985]=25;
cos[11986]=25;
cos[11987]=25;
cos[11988]=25;
cos[11989]=25;
cos[11990]=25;
cos[11991]=25;
cos[11992]=25;
cos[11993]=24;
cos[11994]=24;
cos[11995]=24;
cos[11996]=24;
cos[11997]=24;
cos[11998]=24;
cos[11999]=24;
cos[12000]=24;
cos[12001]=24;
cos[12002]=24;
cos[12003]=24;
cos[12004]=24;
cos[12005]=24;
cos[12006]=24;
cos[12007]=24;
cos[12008]=24;
cos[12009]=24;
cos[12010]=24;
cos[12011]=24;
cos[12012]=24;
cos[12013]=24;
cos[12014]=23;
cos[12015]=23;
cos[12016]=23;
cos[12017]=23;
cos[12018]=23;
cos[12019]=23;
cos[12020]=23;
cos[12021]=23;
cos[12022]=23;
cos[12023]=23;
cos[12024]=23;
cos[12025]=23;
cos[12026]=23;
cos[12027]=23;
cos[12028]=23;
cos[12029]=23;
cos[12030]=23;
cos[12031]=23;
cos[12032]=23;
cos[12033]=23;
cos[12034]=23;
cos[12035]=23;
cos[12036]=22;
cos[12037]=22;
cos[12038]=22;
cos[12039]=22;
cos[12040]=22;
cos[12041]=22;
cos[12042]=22;
cos[12043]=22;
cos[12044]=22;
cos[12045]=22;
cos[12046]=22;
cos[12047]=22;
cos[12048]=22;
cos[12049]=22;
cos[12050]=22;
cos[12051]=22;
cos[12052]=22;
cos[12053]=22;
cos[12054]=22;
cos[12055]=22;
cos[12056]=22;
cos[12057]=21;
cos[12058]=21;
cos[12059]=21;
cos[12060]=21;
cos[12061]=21;
cos[12062]=21;
cos[12063]=21;
cos[12064]=21;
cos[12065]=21;
cos[12066]=21;
cos[12067]=21;
cos[12068]=21;
cos[12069]=21;
cos[12070]=21;
cos[12071]=21;
cos[12072]=21;
cos[12073]=21;
cos[12074]=21;
cos[12075]=21;
cos[12076]=21;
cos[12077]=21;
cos[12078]=20;
cos[12079]=20;
cos[12080]=20;
cos[12081]=20;
cos[12082]=20;
cos[12083]=20;
cos[12084]=20;
cos[12085]=20;
cos[12086]=20;
cos[12087]=20;
cos[12088]=20;
cos[12089]=20;
cos[12090]=20;
cos[12091]=20;
cos[12092]=20;
cos[12093]=20;
cos[12094]=20;
cos[12095]=20;
cos[12096]=20;
cos[12097]=20;
cos[12098]=20;
cos[12099]=19;
cos[12100]=19;
cos[12101]=19;
cos[12102]=19;
cos[12103]=19;
cos[12104]=19;
cos[12105]=19;
cos[12106]=19;
cos[12107]=19;
cos[12108]=19;
cos[12109]=19;
cos[12110]=19;
cos[12111]=19;
cos[12112]=19;
cos[12113]=19;
cos[12114]=19;
cos[12115]=19;
cos[12116]=19;
cos[12117]=19;
cos[12118]=19;
cos[12119]=19;
cos[12120]=18;
cos[12121]=18;
cos[12122]=18;
cos[12123]=18;
cos[12124]=18;
cos[12125]=18;
cos[12126]=18;
cos[12127]=18;
cos[12128]=18;
cos[12129]=18;
cos[12130]=18;
cos[12131]=18;
cos[12132]=18;
cos[12133]=18;
cos[12134]=18;
cos[12135]=18;
cos[12136]=18;
cos[12137]=18;
cos[12138]=18;
cos[12139]=18;
cos[12140]=18;
cos[12141]=17;
cos[12142]=17;
cos[12143]=17;
cos[12144]=17;
cos[12145]=17;
cos[12146]=17;
cos[12147]=17;
cos[12148]=17;
cos[12149]=17;
cos[12150]=17;
cos[12151]=17;
cos[12152]=17;
cos[12153]=17;
cos[12154]=17;
cos[12155]=17;
cos[12156]=17;
cos[12157]=17;
cos[12158]=17;
cos[12159]=17;
cos[12160]=17;
cos[12161]=17;
cos[12162]=16;
cos[12163]=16;
cos[12164]=16;
cos[12165]=16;
cos[12166]=16;
cos[12167]=16;
cos[12168]=16;
cos[12169]=16;
cos[12170]=16;
cos[12171]=16;
cos[12172]=16;
cos[12173]=16;
cos[12174]=16;
cos[12175]=16;
cos[12176]=16;
cos[12177]=16;
cos[12178]=16;
cos[12179]=16;
cos[12180]=16;
cos[12181]=16;
cos[12182]=16;
cos[12183]=15;
cos[12184]=15;
cos[12185]=15;
cos[12186]=15;
cos[12187]=15;
cos[12188]=15;
cos[12189]=15;
cos[12190]=15;
cos[12191]=15;
cos[12192]=15;
cos[12193]=15;
cos[12194]=15;
cos[12195]=15;
cos[12196]=15;
cos[12197]=15;
cos[12198]=15;
cos[12199]=15;
cos[12200]=15;
cos[12201]=15;
cos[12202]=15;
cos[12203]=14;
cos[12204]=14;
cos[12205]=14;
cos[12206]=14;
cos[12207]=14;
cos[12208]=14;
cos[12209]=14;
cos[12210]=14;
cos[12211]=14;
cos[12212]=14;
cos[12213]=14;
cos[12214]=14;
cos[12215]=14;
cos[12216]=14;
cos[12217]=14;
cos[12218]=14;
cos[12219]=14;
cos[12220]=14;
cos[12221]=14;
cos[12222]=14;
cos[12223]=14;
cos[12224]=13;
cos[12225]=13;
cos[12226]=13;
cos[12227]=13;
cos[12228]=13;
cos[12229]=13;
cos[12230]=13;
cos[12231]=13;
cos[12232]=13;
cos[12233]=13;
cos[12234]=13;
cos[12235]=13;
cos[12236]=13;
cos[12237]=13;
cos[12238]=13;
cos[12239]=13;
cos[12240]=13;
cos[12241]=13;
cos[12242]=13;
cos[12243]=13;
cos[12244]=13;
cos[12245]=12;
cos[12246]=12;
cos[12247]=12;
cos[12248]=12;
cos[12249]=12;
cos[12250]=12;
cos[12251]=12;
cos[12252]=12;
cos[12253]=12;
cos[12254]=12;
cos[12255]=12;
cos[12256]=12;
cos[12257]=12;
cos[12258]=12;
cos[12259]=12;
cos[12260]=12;
cos[12261]=12;
cos[12262]=12;
cos[12263]=12;
cos[12264]=12;
cos[12265]=11;
cos[12266]=11;
cos[12267]=11;
cos[12268]=11;
cos[12269]=11;
cos[12270]=11;
cos[12271]=11;
cos[12272]=11;
cos[12273]=11;
cos[12274]=11;
cos[12275]=11;
cos[12276]=11;
cos[12277]=11;
cos[12278]=11;
cos[12279]=11;
cos[12280]=11;
cos[12281]=11;
cos[12282]=11;
cos[12283]=11;
cos[12284]=11;
cos[12285]=11;
cos[12286]=10;
cos[12287]=10;
cos[12288]=10;
cos[12289]=10;
cos[12290]=10;
cos[12291]=10;
cos[12292]=10;
cos[12293]=10;
cos[12294]=10;
cos[12295]=10;
cos[12296]=10;
cos[12297]=10;
cos[12298]=10;
cos[12299]=10;
cos[12300]=10;
cos[12301]=10;
cos[12302]=10;
cos[12303]=10;
cos[12304]=10;
cos[12305]=10;
cos[12306]=9;
cos[12307]=9;
cos[12308]=9;
cos[12309]=9;
cos[12310]=9;
cos[12311]=9;
cos[12312]=9;
cos[12313]=9;
cos[12314]=9;
cos[12315]=9;
cos[12316]=9;
cos[12317]=9;
cos[12318]=9;
cos[12319]=9;
cos[12320]=9;
cos[12321]=9;
cos[12322]=9;
cos[12323]=9;
cos[12324]=9;
cos[12325]=9;
cos[12326]=9;
cos[12327]=8;
cos[12328]=8;
cos[12329]=8;
cos[12330]=8;
cos[12331]=8;
cos[12332]=8;
cos[12333]=8;
cos[12334]=8;
cos[12335]=8;
cos[12336]=8;
cos[12337]=8;
cos[12338]=8;
cos[12339]=8;
cos[12340]=8;
cos[12341]=8;
cos[12342]=8;
cos[12343]=8;
cos[12344]=8;
cos[12345]=8;
cos[12346]=8;
cos[12347]=7;
cos[12348]=7;
cos[12349]=7;
cos[12350]=7;
cos[12351]=7;
cos[12352]=7;
cos[12353]=7;
cos[12354]=7;
cos[12355]=7;
cos[12356]=7;
cos[12357]=7;
cos[12358]=7;
cos[12359]=7;
cos[12360]=7;
cos[12361]=7;
cos[12362]=7;
cos[12363]=7;
cos[12364]=7;
cos[12365]=7;
cos[12366]=7;
cos[12367]=7;
cos[12368]=6;
cos[12369]=6;
cos[12370]=6;
cos[12371]=6;
cos[12372]=6;
cos[12373]=6;
cos[12374]=6;
cos[12375]=6;
cos[12376]=6;
cos[12377]=6;
cos[12378]=6;
cos[12379]=6;
cos[12380]=6;
cos[12381]=6;
cos[12382]=6;
cos[12383]=6;
cos[12384]=6;
cos[12385]=6;
cos[12386]=6;
cos[12387]=6;
cos[12388]=5;
cos[12389]=5;
cos[12390]=5;
cos[12391]=5;
cos[12392]=5;
cos[12393]=5;
cos[12394]=5;
cos[12395]=5;
cos[12396]=5;
cos[12397]=5;
cos[12398]=5;
cos[12399]=5;
cos[12400]=5;
cos[12401]=5;
cos[12402]=5;
cos[12403]=5;
cos[12404]=5;
cos[12405]=5;
cos[12406]=5;
cos[12407]=5;
cos[12408]=5;
cos[12409]=4;
cos[12410]=4;
cos[12411]=4;
cos[12412]=4;
cos[12413]=4;
cos[12414]=4;
cos[12415]=4;
cos[12416]=4;
cos[12417]=4;
cos[12418]=4;
cos[12419]=4;
cos[12420]=4;
cos[12421]=4;
cos[12422]=4;
cos[12423]=4;
cos[12424]=4;
cos[12425]=4;
cos[12426]=4;
cos[12427]=4;
cos[12428]=4;
cos[12429]=3;
cos[12430]=3;
cos[12431]=3;
cos[12432]=3;
cos[12433]=3;
cos[12434]=3;
cos[12435]=3;
cos[12436]=3;
cos[12437]=3;
cos[12438]=3;
cos[12439]=3;
cos[12440]=3;
cos[12441]=3;
cos[12442]=3;
cos[12443]=3;
cos[12444]=3;
cos[12445]=3;
cos[12446]=3;
cos[12447]=3;
cos[12448]=3;
cos[12449]=3;
cos[12450]=2;
cos[12451]=2;
cos[12452]=2;
cos[12453]=2;
cos[12454]=2;
cos[12455]=2;
cos[12456]=2;
cos[12457]=2;
cos[12458]=2;
cos[12459]=2;
cos[12460]=2;
cos[12461]=2;
cos[12462]=2;
cos[12463]=2;
cos[12464]=2;
cos[12465]=2;
cos[12466]=2;
cos[12467]=2;
cos[12468]=2;
cos[12469]=2;
cos[12470]=1;
cos[12471]=1;
cos[12472]=1;
cos[12473]=1;
cos[12474]=1;
cos[12475]=1;
cos[12476]=1;
cos[12477]=1;
cos[12478]=1;
cos[12479]=1;
cos[12480]=1;
cos[12481]=1;
cos[12482]=1;
cos[12483]=1;
cos[12484]=1;
cos[12485]=1;
cos[12486]=1;
cos[12487]=1;
cos[12488]=1;
cos[12489]=1;
cos[12490]=0;
cos[12491]=0;
cos[12492]=0;
cos[12493]=0;
cos[12494]=0;
cos[12495]=0;
cos[12496]=0;
cos[12497]=0;
cos[12498]=0;
cos[12499]=0;
cos[12500]=0;
cos[12501]=0;
cos[12502]=0;
cos[12503]=0;
cos[12504]=0;
cos[12505]=0;
cos[12506]=0;
cos[12507]=0;
cos[12508]=0;
cos[12509]=0;
cos[12510]=0;
cos[12511]=-1;
cos[12512]=-1;
cos[12513]=-1;
cos[12514]=-1;
cos[12515]=-1;
cos[12516]=-1;
cos[12517]=-1;
cos[12518]=-1;
cos[12519]=-1;
cos[12520]=-1;
cos[12521]=-1;
cos[12522]=-1;
cos[12523]=-1;
cos[12524]=-1;
cos[12525]=-1;
cos[12526]=-1;
cos[12527]=-1;
cos[12528]=-1;
cos[12529]=-1;
cos[12530]=-1;
cos[12531]=-2;
cos[12532]=-2;
cos[12533]=-2;
cos[12534]=-2;
cos[12535]=-2;
cos[12536]=-2;
cos[12537]=-2;
cos[12538]=-2;
cos[12539]=-2;
cos[12540]=-2;
cos[12541]=-2;
cos[12542]=-2;
cos[12543]=-2;
cos[12544]=-2;
cos[12545]=-2;
cos[12546]=-2;
cos[12547]=-2;
cos[12548]=-2;
cos[12549]=-2;
cos[12550]=-2;
cos[12551]=-3;
cos[12552]=-3;
cos[12553]=-3;
cos[12554]=-3;
cos[12555]=-3;
cos[12556]=-3;
cos[12557]=-3;
cos[12558]=-3;
cos[12559]=-3;
cos[12560]=-3;
cos[12561]=-3;
cos[12562]=-3;
cos[12563]=-3;
cos[12564]=-3;
cos[12565]=-3;
cos[12566]=-3;
cos[12567]=-3;
cos[12568]=-3;
cos[12569]=-3;
cos[12570]=-3;
cos[12571]=-3;
cos[12572]=-4;
cos[12573]=-4;
cos[12574]=-4;
cos[12575]=-4;
cos[12576]=-4;
cos[12577]=-4;
cos[12578]=-4;
cos[12579]=-4;
cos[12580]=-4;
cos[12581]=-4;
cos[12582]=-4;
cos[12583]=-4;
cos[12584]=-4;
cos[12585]=-4;
cos[12586]=-4;
cos[12587]=-4;
cos[12588]=-4;
cos[12589]=-4;
cos[12590]=-4;
cos[12591]=-4;
cos[12592]=-5;
cos[12593]=-5;
cos[12594]=-5;
cos[12595]=-5;
cos[12596]=-5;
cos[12597]=-5;
cos[12598]=-5;
cos[12599]=-5;
cos[12600]=-5;
cos[12601]=-5;
cos[12602]=-5;
cos[12603]=-5;
cos[12604]=-5;
cos[12605]=-5;
cos[12606]=-5;
cos[12607]=-5;
cos[12608]=-5;
cos[12609]=-5;
cos[12610]=-5;
cos[12611]=-5;
cos[12612]=-5;
cos[12613]=-6;
cos[12614]=-6;
cos[12615]=-6;
cos[12616]=-6;
cos[12617]=-6;
cos[12618]=-6;
cos[12619]=-6;
cos[12620]=-6;
cos[12621]=-6;
cos[12622]=-6;
cos[12623]=-6;
cos[12624]=-6;
cos[12625]=-6;
cos[12626]=-6;
cos[12627]=-6;
cos[12628]=-6;
cos[12629]=-6;
cos[12630]=-6;
cos[12631]=-6;
cos[12632]=-6;
cos[12633]=-7;
cos[12634]=-7;
cos[12635]=-7;
cos[12636]=-7;
cos[12637]=-7;
cos[12638]=-7;
cos[12639]=-7;
cos[12640]=-7;
cos[12641]=-7;
cos[12642]=-7;
cos[12643]=-7;
cos[12644]=-7;
cos[12645]=-7;
cos[12646]=-7;
cos[12647]=-7;
cos[12648]=-7;
cos[12649]=-7;
cos[12650]=-7;
cos[12651]=-7;
cos[12652]=-7;
cos[12653]=-7;
cos[12654]=-8;
cos[12655]=-8;
cos[12656]=-8;
cos[12657]=-8;
cos[12658]=-8;
cos[12659]=-8;
cos[12660]=-8;
cos[12661]=-8;
cos[12662]=-8;
cos[12663]=-8;
cos[12664]=-8;
cos[12665]=-8;
cos[12666]=-8;
cos[12667]=-8;
cos[12668]=-8;
cos[12669]=-8;
cos[12670]=-8;
cos[12671]=-8;
cos[12672]=-8;
cos[12673]=-8;
cos[12674]=-9;
cos[12675]=-9;
cos[12676]=-9;
cos[12677]=-9;
cos[12678]=-9;
cos[12679]=-9;
cos[12680]=-9;
cos[12681]=-9;
cos[12682]=-9;
cos[12683]=-9;
cos[12684]=-9;
cos[12685]=-9;
cos[12686]=-9;
cos[12687]=-9;
cos[12688]=-9;
cos[12689]=-9;
cos[12690]=-9;
cos[12691]=-9;
cos[12692]=-9;
cos[12693]=-9;
cos[12694]=-9;
cos[12695]=-10;
cos[12696]=-10;
cos[12697]=-10;
cos[12698]=-10;
cos[12699]=-10;
cos[12700]=-10;
cos[12701]=-10;
cos[12702]=-10;
cos[12703]=-10;
cos[12704]=-10;
cos[12705]=-10;
cos[12706]=-10;
cos[12707]=-10;
cos[12708]=-10;
cos[12709]=-10;
cos[12710]=-10;
cos[12711]=-10;
cos[12712]=-10;
cos[12713]=-10;
cos[12714]=-10;
cos[12715]=-11;
cos[12716]=-11;
cos[12717]=-11;
cos[12718]=-11;
cos[12719]=-11;
cos[12720]=-11;
cos[12721]=-11;
cos[12722]=-11;
cos[12723]=-11;
cos[12724]=-11;
cos[12725]=-11;
cos[12726]=-11;
cos[12727]=-11;
cos[12728]=-11;
cos[12729]=-11;
cos[12730]=-11;
cos[12731]=-11;
cos[12732]=-11;
cos[12733]=-11;
cos[12734]=-11;
cos[12735]=-11;
cos[12736]=-12;
cos[12737]=-12;
cos[12738]=-12;
cos[12739]=-12;
cos[12740]=-12;
cos[12741]=-12;
cos[12742]=-12;
cos[12743]=-12;
cos[12744]=-12;
cos[12745]=-12;
cos[12746]=-12;
cos[12747]=-12;
cos[12748]=-12;
cos[12749]=-12;
cos[12750]=-12;
cos[12751]=-12;
cos[12752]=-12;
cos[12753]=-12;
cos[12754]=-12;
cos[12755]=-12;
cos[12756]=-13;
cos[12757]=-13;
cos[12758]=-13;
cos[12759]=-13;
cos[12760]=-13;
cos[12761]=-13;
cos[12762]=-13;
cos[12763]=-13;
cos[12764]=-13;
cos[12765]=-13;
cos[12766]=-13;
cos[12767]=-13;
cos[12768]=-13;
cos[12769]=-13;
cos[12770]=-13;
cos[12771]=-13;
cos[12772]=-13;
cos[12773]=-13;
cos[12774]=-13;
cos[12775]=-13;
cos[12776]=-13;
cos[12777]=-14;
cos[12778]=-14;
cos[12779]=-14;
cos[12780]=-14;
cos[12781]=-14;
cos[12782]=-14;
cos[12783]=-14;
cos[12784]=-14;
cos[12785]=-14;
cos[12786]=-14;
cos[12787]=-14;
cos[12788]=-14;
cos[12789]=-14;
cos[12790]=-14;
cos[12791]=-14;
cos[12792]=-14;
cos[12793]=-14;
cos[12794]=-14;
cos[12795]=-14;
cos[12796]=-14;
cos[12797]=-14;
cos[12798]=-15;
cos[12799]=-15;
cos[12800]=-15;
cos[12801]=-15;
cos[12802]=-15;
cos[12803]=-15;
cos[12804]=-15;
cos[12805]=-15;
cos[12806]=-15;
cos[12807]=-15;
cos[12808]=-15;
cos[12809]=-15;
cos[12810]=-15;
cos[12811]=-15;
cos[12812]=-15;
cos[12813]=-15;
cos[12814]=-15;
cos[12815]=-15;
cos[12816]=-15;
cos[12817]=-15;
cos[12818]=-16;
cos[12819]=-16;
cos[12820]=-16;
cos[12821]=-16;
cos[12822]=-16;
cos[12823]=-16;
cos[12824]=-16;
cos[12825]=-16;
cos[12826]=-16;
cos[12827]=-16;
cos[12828]=-16;
cos[12829]=-16;
cos[12830]=-16;
cos[12831]=-16;
cos[12832]=-16;
cos[12833]=-16;
cos[12834]=-16;
cos[12835]=-16;
cos[12836]=-16;
cos[12837]=-16;
cos[12838]=-16;
cos[12839]=-17;
cos[12840]=-17;
cos[12841]=-17;
cos[12842]=-17;
cos[12843]=-17;
cos[12844]=-17;
cos[12845]=-17;
cos[12846]=-17;
cos[12847]=-17;
cos[12848]=-17;
cos[12849]=-17;
cos[12850]=-17;
cos[12851]=-17;
cos[12852]=-17;
cos[12853]=-17;
cos[12854]=-17;
cos[12855]=-17;
cos[12856]=-17;
cos[12857]=-17;
cos[12858]=-17;
cos[12859]=-17;
cos[12860]=-18;
cos[12861]=-18;
cos[12862]=-18;
cos[12863]=-18;
cos[12864]=-18;
cos[12865]=-18;
cos[12866]=-18;
cos[12867]=-18;
cos[12868]=-18;
cos[12869]=-18;
cos[12870]=-18;
cos[12871]=-18;
cos[12872]=-18;
cos[12873]=-18;
cos[12874]=-18;
cos[12875]=-18;
cos[12876]=-18;
cos[12877]=-18;
cos[12878]=-18;
cos[12879]=-18;
cos[12880]=-18;
cos[12881]=-19;
cos[12882]=-19;
cos[12883]=-19;
cos[12884]=-19;
cos[12885]=-19;
cos[12886]=-19;
cos[12887]=-19;
cos[12888]=-19;
cos[12889]=-19;
cos[12890]=-19;
cos[12891]=-19;
cos[12892]=-19;
cos[12893]=-19;
cos[12894]=-19;
cos[12895]=-19;
cos[12896]=-19;
cos[12897]=-19;
cos[12898]=-19;
cos[12899]=-19;
cos[12900]=-19;
cos[12901]=-19;
cos[12902]=-20;
cos[12903]=-20;
cos[12904]=-20;
cos[12905]=-20;
cos[12906]=-20;
cos[12907]=-20;
cos[12908]=-20;
cos[12909]=-20;
cos[12910]=-20;
cos[12911]=-20;
cos[12912]=-20;
cos[12913]=-20;
cos[12914]=-20;
cos[12915]=-20;
cos[12916]=-20;
cos[12917]=-20;
cos[12918]=-20;
cos[12919]=-20;
cos[12920]=-20;
cos[12921]=-20;
cos[12922]=-20;
cos[12923]=-21;
cos[12924]=-21;
cos[12925]=-21;
cos[12926]=-21;
cos[12927]=-21;
cos[12928]=-21;
cos[12929]=-21;
cos[12930]=-21;
cos[12931]=-21;
cos[12932]=-21;
cos[12933]=-21;
cos[12934]=-21;
cos[12935]=-21;
cos[12936]=-21;
cos[12937]=-21;
cos[12938]=-21;
cos[12939]=-21;
cos[12940]=-21;
cos[12941]=-21;
cos[12942]=-21;
cos[12943]=-21;
cos[12944]=-22;
cos[12945]=-22;
cos[12946]=-22;
cos[12947]=-22;
cos[12948]=-22;
cos[12949]=-22;
cos[12950]=-22;
cos[12951]=-22;
cos[12952]=-22;
cos[12953]=-22;
cos[12954]=-22;
cos[12955]=-22;
cos[12956]=-22;
cos[12957]=-22;
cos[12958]=-22;
cos[12959]=-22;
cos[12960]=-22;
cos[12961]=-22;
cos[12962]=-22;
cos[12963]=-22;
cos[12964]=-22;
cos[12965]=-23;
cos[12966]=-23;
cos[12967]=-23;
cos[12968]=-23;
cos[12969]=-23;
cos[12970]=-23;
cos[12971]=-23;
cos[12972]=-23;
cos[12973]=-23;
cos[12974]=-23;
cos[12975]=-23;
cos[12976]=-23;
cos[12977]=-23;
cos[12978]=-23;
cos[12979]=-23;
cos[12980]=-23;
cos[12981]=-23;
cos[12982]=-23;
cos[12983]=-23;
cos[12984]=-23;
cos[12985]=-23;
cos[12986]=-23;
cos[12987]=-24;
cos[12988]=-24;
cos[12989]=-24;
cos[12990]=-24;
cos[12991]=-24;
cos[12992]=-24;
cos[12993]=-24;
cos[12994]=-24;
cos[12995]=-24;
cos[12996]=-24;
cos[12997]=-24;
cos[12998]=-24;
cos[12999]=-24;
cos[13000]=-24;
cos[13001]=-24;
cos[13002]=-24;
cos[13003]=-24;
cos[13004]=-24;
cos[13005]=-24;
cos[13006]=-24;
cos[13007]=-24;
cos[13008]=-25;
cos[13009]=-25;
cos[13010]=-25;
cos[13011]=-25;
cos[13012]=-25;
cos[13013]=-25;
cos[13014]=-25;
cos[13015]=-25;
cos[13016]=-25;
cos[13017]=-25;
cos[13018]=-25;
cos[13019]=-25;
cos[13020]=-25;
cos[13021]=-25;
cos[13022]=-25;
cos[13023]=-25;
cos[13024]=-25;
cos[13025]=-25;
cos[13026]=-25;
cos[13027]=-25;
cos[13028]=-25;
cos[13029]=-25;
cos[13030]=-26;
cos[13031]=-26;
cos[13032]=-26;
cos[13033]=-26;
cos[13034]=-26;
cos[13035]=-26;
cos[13036]=-26;
cos[13037]=-26;
cos[13038]=-26;
cos[13039]=-26;
cos[13040]=-26;
cos[13041]=-26;
cos[13042]=-26;
cos[13043]=-26;
cos[13044]=-26;
cos[13045]=-26;
cos[13046]=-26;
cos[13047]=-26;
cos[13048]=-26;
cos[13049]=-26;
cos[13050]=-26;
cos[13051]=-27;
cos[13052]=-27;
cos[13053]=-27;
cos[13054]=-27;
cos[13055]=-27;
cos[13056]=-27;
cos[13057]=-27;
cos[13058]=-27;
cos[13059]=-27;
cos[13060]=-27;
cos[13061]=-27;
cos[13062]=-27;
cos[13063]=-27;
cos[13064]=-27;
cos[13065]=-27;
cos[13066]=-27;
cos[13067]=-27;
cos[13068]=-27;
cos[13069]=-27;
cos[13070]=-27;
cos[13071]=-27;
cos[13072]=-27;
cos[13073]=-28;
cos[13074]=-28;
cos[13075]=-28;
cos[13076]=-28;
cos[13077]=-28;
cos[13078]=-28;
cos[13079]=-28;
cos[13080]=-28;
cos[13081]=-28;
cos[13082]=-28;
cos[13083]=-28;
cos[13084]=-28;
cos[13085]=-28;
cos[13086]=-28;
cos[13087]=-28;
cos[13088]=-28;
cos[13089]=-28;
cos[13090]=-28;
cos[13091]=-28;
cos[13092]=-28;
cos[13093]=-28;
cos[13094]=-28;
cos[13095]=-29;
cos[13096]=-29;
cos[13097]=-29;
cos[13098]=-29;
cos[13099]=-29;
cos[13100]=-29;
cos[13101]=-29;
cos[13102]=-29;
cos[13103]=-29;
cos[13104]=-29;
cos[13105]=-29;
cos[13106]=-29;
cos[13107]=-29;
cos[13108]=-29;
cos[13109]=-29;
cos[13110]=-29;
cos[13111]=-29;
cos[13112]=-29;
cos[13113]=-29;
cos[13114]=-29;
cos[13115]=-29;
cos[13116]=-29;
cos[13117]=-30;
cos[13118]=-30;
cos[13119]=-30;
cos[13120]=-30;
cos[13121]=-30;
cos[13122]=-30;
cos[13123]=-30;
cos[13124]=-30;
cos[13125]=-30;
cos[13126]=-30;
cos[13127]=-30;
cos[13128]=-30;
cos[13129]=-30;
cos[13130]=-30;
cos[13131]=-30;
cos[13132]=-30;
cos[13133]=-30;
cos[13134]=-30;
cos[13135]=-30;
cos[13136]=-30;
cos[13137]=-30;
cos[13138]=-30;
cos[13139]=-31;
cos[13140]=-31;
cos[13141]=-31;
cos[13142]=-31;
cos[13143]=-31;
cos[13144]=-31;
cos[13145]=-31;
cos[13146]=-31;
cos[13147]=-31;
cos[13148]=-31;
cos[13149]=-31;
cos[13150]=-31;
cos[13151]=-31;
cos[13152]=-31;
cos[13153]=-31;
cos[13154]=-31;
cos[13155]=-31;
cos[13156]=-31;
cos[13157]=-31;
cos[13158]=-31;
cos[13159]=-31;
cos[13160]=-31;
cos[13161]=-32;
cos[13162]=-32;
cos[13163]=-32;
cos[13164]=-32;
cos[13165]=-32;
cos[13166]=-32;
cos[13167]=-32;
cos[13168]=-32;
cos[13169]=-32;
cos[13170]=-32;
cos[13171]=-32;
cos[13172]=-32;
cos[13173]=-32;
cos[13174]=-32;
cos[13175]=-32;
cos[13176]=-32;
cos[13177]=-32;
cos[13178]=-32;
cos[13179]=-32;
cos[13180]=-32;
cos[13181]=-32;
cos[13182]=-32;
cos[13183]=-33;
cos[13184]=-33;
cos[13185]=-33;
cos[13186]=-33;
cos[13187]=-33;
cos[13188]=-33;
cos[13189]=-33;
cos[13190]=-33;
cos[13191]=-33;
cos[13192]=-33;
cos[13193]=-33;
cos[13194]=-33;
cos[13195]=-33;
cos[13196]=-33;
cos[13197]=-33;
cos[13198]=-33;
cos[13199]=-33;
cos[13200]=-33;
cos[13201]=-33;
cos[13202]=-33;
cos[13203]=-33;
cos[13204]=-33;
cos[13205]=-33;
cos[13206]=-34;
cos[13207]=-34;
cos[13208]=-34;
cos[13209]=-34;
cos[13210]=-34;
cos[13211]=-34;
cos[13212]=-34;
cos[13213]=-34;
cos[13214]=-34;
cos[13215]=-34;
cos[13216]=-34;
cos[13217]=-34;
cos[13218]=-34;
cos[13219]=-34;
cos[13220]=-34;
cos[13221]=-34;
cos[13222]=-34;
cos[13223]=-34;
cos[13224]=-34;
cos[13225]=-34;
cos[13226]=-34;
cos[13227]=-34;
cos[13228]=-35;
cos[13229]=-35;
cos[13230]=-35;
cos[13231]=-35;
cos[13232]=-35;
cos[13233]=-35;
cos[13234]=-35;
cos[13235]=-35;
cos[13236]=-35;
cos[13237]=-35;
cos[13238]=-35;
cos[13239]=-35;
cos[13240]=-35;
cos[13241]=-35;
cos[13242]=-35;
cos[13243]=-35;
cos[13244]=-35;
cos[13245]=-35;
cos[13246]=-35;
cos[13247]=-35;
cos[13248]=-35;
cos[13249]=-35;
cos[13250]=-35;
cos[13251]=-36;
cos[13252]=-36;
cos[13253]=-36;
cos[13254]=-36;
cos[13255]=-36;
cos[13256]=-36;
cos[13257]=-36;
cos[13258]=-36;
cos[13259]=-36;
cos[13260]=-36;
cos[13261]=-36;
cos[13262]=-36;
cos[13263]=-36;
cos[13264]=-36;
cos[13265]=-36;
cos[13266]=-36;
cos[13267]=-36;
cos[13268]=-36;
cos[13269]=-36;
cos[13270]=-36;
cos[13271]=-36;
cos[13272]=-36;
cos[13273]=-36;
cos[13274]=-37;
cos[13275]=-37;
cos[13276]=-37;
cos[13277]=-37;
cos[13278]=-37;
cos[13279]=-37;
cos[13280]=-37;
cos[13281]=-37;
cos[13282]=-37;
cos[13283]=-37;
cos[13284]=-37;
cos[13285]=-37;
cos[13286]=-37;
cos[13287]=-37;
cos[13288]=-37;
cos[13289]=-37;
cos[13290]=-37;
cos[13291]=-37;
cos[13292]=-37;
cos[13293]=-37;
cos[13294]=-37;
cos[13295]=-37;
cos[13296]=-37;
cos[13297]=-38;
cos[13298]=-38;
cos[13299]=-38;
cos[13300]=-38;
cos[13301]=-38;
cos[13302]=-38;
cos[13303]=-38;
cos[13304]=-38;
cos[13305]=-38;
cos[13306]=-38;
cos[13307]=-38;
cos[13308]=-38;
cos[13309]=-38;
cos[13310]=-38;
cos[13311]=-38;
cos[13312]=-38;
cos[13313]=-38;
cos[13314]=-38;
cos[13315]=-38;
cos[13316]=-38;
cos[13317]=-38;
cos[13318]=-38;
cos[13319]=-38;
cos[13320]=-38;
cos[13321]=-39;
cos[13322]=-39;
cos[13323]=-39;
cos[13324]=-39;
cos[13325]=-39;
cos[13326]=-39;
cos[13327]=-39;
cos[13328]=-39;
cos[13329]=-39;
cos[13330]=-39;
cos[13331]=-39;
cos[13332]=-39;
cos[13333]=-39;
cos[13334]=-39;
cos[13335]=-39;
cos[13336]=-39;
cos[13337]=-39;
cos[13338]=-39;
cos[13339]=-39;
cos[13340]=-39;
cos[13341]=-39;
cos[13342]=-39;
cos[13343]=-39;
cos[13344]=-40;
cos[13345]=-40;
cos[13346]=-40;
cos[13347]=-40;
cos[13348]=-40;
cos[13349]=-40;
cos[13350]=-40;
cos[13351]=-40;
cos[13352]=-40;
cos[13353]=-40;
cos[13354]=-40;
cos[13355]=-40;
cos[13356]=-40;
cos[13357]=-40;
cos[13358]=-40;
cos[13359]=-40;
cos[13360]=-40;
cos[13361]=-40;
cos[13362]=-40;
cos[13363]=-40;
cos[13364]=-40;
cos[13365]=-40;
cos[13366]=-40;
cos[13367]=-40;
cos[13368]=-41;
cos[13369]=-41;
cos[13370]=-41;
cos[13371]=-41;
cos[13372]=-41;
cos[13373]=-41;
cos[13374]=-41;
cos[13375]=-41;
cos[13376]=-41;
cos[13377]=-41;
cos[13378]=-41;
cos[13379]=-41;
cos[13380]=-41;
cos[13381]=-41;
cos[13382]=-41;
cos[13383]=-41;
cos[13384]=-41;
cos[13385]=-41;
cos[13386]=-41;
cos[13387]=-41;
cos[13388]=-41;
cos[13389]=-41;
cos[13390]=-41;
cos[13391]=-41;
cos[13392]=-42;
cos[13393]=-42;
cos[13394]=-42;
cos[13395]=-42;
cos[13396]=-42;
cos[13397]=-42;
cos[13398]=-42;
cos[13399]=-42;
cos[13400]=-42;
cos[13401]=-42;
cos[13402]=-42;
cos[13403]=-42;
cos[13404]=-42;
cos[13405]=-42;
cos[13406]=-42;
cos[13407]=-42;
cos[13408]=-42;
cos[13409]=-42;
cos[13410]=-42;
cos[13411]=-42;
cos[13412]=-42;
cos[13413]=-42;
cos[13414]=-42;
cos[13415]=-42;
cos[13416]=-43;
cos[13417]=-43;
cos[13418]=-43;
cos[13419]=-43;
cos[13420]=-43;
cos[13421]=-43;
cos[13422]=-43;
cos[13423]=-43;
cos[13424]=-43;
cos[13425]=-43;
cos[13426]=-43;
cos[13427]=-43;
cos[13428]=-43;
cos[13429]=-43;
cos[13430]=-43;
cos[13431]=-43;
cos[13432]=-43;
cos[13433]=-43;
cos[13434]=-43;
cos[13435]=-43;
cos[13436]=-43;
cos[13437]=-43;
cos[13438]=-43;
cos[13439]=-43;
cos[13440]=-44;
cos[13441]=-44;
cos[13442]=-44;
cos[13443]=-44;
cos[13444]=-44;
cos[13445]=-44;
cos[13446]=-44;
cos[13447]=-44;
cos[13448]=-44;
cos[13449]=-44;
cos[13450]=-44;
cos[13451]=-44;
cos[13452]=-44;
cos[13453]=-44;
cos[13454]=-44;
cos[13455]=-44;
cos[13456]=-44;
cos[13457]=-44;
cos[13458]=-44;
cos[13459]=-44;
cos[13460]=-44;
cos[13461]=-44;
cos[13462]=-44;
cos[13463]=-44;
cos[13464]=-44;
cos[13465]=-45;
cos[13466]=-45;
cos[13467]=-45;
cos[13468]=-45;
cos[13469]=-45;
cos[13470]=-45;
cos[13471]=-45;
cos[13472]=-45;
cos[13473]=-45;
cos[13474]=-45;
cos[13475]=-45;
cos[13476]=-45;
cos[13477]=-45;
cos[13478]=-45;
cos[13479]=-45;
cos[13480]=-45;
cos[13481]=-45;
cos[13482]=-45;
cos[13483]=-45;
cos[13484]=-45;
cos[13485]=-45;
cos[13486]=-45;
cos[13487]=-45;
cos[13488]=-45;
cos[13489]=-45;
cos[13490]=-46;
cos[13491]=-46;
cos[13492]=-46;
cos[13493]=-46;
cos[13494]=-46;
cos[13495]=-46;
cos[13496]=-46;
cos[13497]=-46;
cos[13498]=-46;
cos[13499]=-46;
cos[13500]=-46;
cos[13501]=-46;
cos[13502]=-46;
cos[13503]=-46;
cos[13504]=-46;
cos[13505]=-46;
cos[13506]=-46;
cos[13507]=-46;
cos[13508]=-46;
cos[13509]=-46;
cos[13510]=-46;
cos[13511]=-46;
cos[13512]=-46;
cos[13513]=-46;
cos[13514]=-46;
cos[13515]=-47;
cos[13516]=-47;
cos[13517]=-47;
cos[13518]=-47;
cos[13519]=-47;
cos[13520]=-47;
cos[13521]=-47;
cos[13522]=-47;
cos[13523]=-47;
cos[13524]=-47;
cos[13525]=-47;
cos[13526]=-47;
cos[13527]=-47;
cos[13528]=-47;
cos[13529]=-47;
cos[13530]=-47;
cos[13531]=-47;
cos[13532]=-47;
cos[13533]=-47;
cos[13534]=-47;
cos[13535]=-47;
cos[13536]=-47;
cos[13537]=-47;
cos[13538]=-47;
cos[13539]=-47;
cos[13540]=-47;
cos[13541]=-48;
cos[13542]=-48;
cos[13543]=-48;
cos[13544]=-48;
cos[13545]=-48;
cos[13546]=-48;
cos[13547]=-48;
cos[13548]=-48;
cos[13549]=-48;
cos[13550]=-48;
cos[13551]=-48;
cos[13552]=-48;
cos[13553]=-48;
cos[13554]=-48;
cos[13555]=-48;
cos[13556]=-48;
cos[13557]=-48;
cos[13558]=-48;
cos[13559]=-48;
cos[13560]=-48;
cos[13561]=-48;
cos[13562]=-48;
cos[13563]=-48;
cos[13564]=-48;
cos[13565]=-48;
cos[13566]=-49;
cos[13567]=-49;
cos[13568]=-49;
cos[13569]=-49;
cos[13570]=-49;
cos[13571]=-49;
cos[13572]=-49;
cos[13573]=-49;
cos[13574]=-49;
cos[13575]=-49;
cos[13576]=-49;
cos[13577]=-49;
cos[13578]=-49;
cos[13579]=-49;
cos[13580]=-49;
cos[13581]=-49;
cos[13582]=-49;
cos[13583]=-49;
cos[13584]=-49;
cos[13585]=-49;
cos[13586]=-49;
cos[13587]=-49;
cos[13588]=-49;
cos[13589]=-49;
cos[13590]=-49;
cos[13591]=-49;
cos[13592]=-49;
cos[13593]=-50;
cos[13594]=-50;
cos[13595]=-50;
cos[13596]=-50;
cos[13597]=-50;
cos[13598]=-50;
cos[13599]=-50;
cos[13600]=-50;
cos[13601]=-50;
cos[13602]=-50;
cos[13603]=-50;
cos[13604]=-50;
cos[13605]=-50;
cos[13606]=-50;
cos[13607]=-50;
cos[13608]=-50;
cos[13609]=-50;
cos[13610]=-50;
cos[13611]=-50;
cos[13612]=-50;
cos[13613]=-50;
cos[13614]=-50;
cos[13615]=-50;
cos[13616]=-50;
cos[13617]=-50;
cos[13618]=-50;
cos[13619]=-51;
cos[13620]=-51;
cos[13621]=-51;
cos[13622]=-51;
cos[13623]=-51;
cos[13624]=-51;
cos[13625]=-51;
cos[13626]=-51;
cos[13627]=-51;
cos[13628]=-51;
cos[13629]=-51;
cos[13630]=-51;
cos[13631]=-51;
cos[13632]=-51;
cos[13633]=-51;
cos[13634]=-51;
cos[13635]=-51;
cos[13636]=-51;
cos[13637]=-51;
cos[13638]=-51;
cos[13639]=-51;
cos[13640]=-51;
cos[13641]=-51;
cos[13642]=-51;
cos[13643]=-51;
cos[13644]=-51;
cos[13645]=-51;
cos[13646]=-52;
cos[13647]=-52;
cos[13648]=-52;
cos[13649]=-52;
cos[13650]=-52;
cos[13651]=-52;
cos[13652]=-52;
cos[13653]=-52;
cos[13654]=-52;
cos[13655]=-52;
cos[13656]=-52;
cos[13657]=-52;
cos[13658]=-52;
cos[13659]=-52;
cos[13660]=-52;
cos[13661]=-52;
cos[13662]=-52;
cos[13663]=-52;
cos[13664]=-52;
cos[13665]=-52;
cos[13666]=-52;
cos[13667]=-52;
cos[13668]=-52;
cos[13669]=-52;
cos[13670]=-52;
cos[13671]=-52;
cos[13672]=-52;
cos[13673]=-53;
cos[13674]=-53;
cos[13675]=-53;
cos[13676]=-53;
cos[13677]=-53;
cos[13678]=-53;
cos[13679]=-53;
cos[13680]=-53;
cos[13681]=-53;
cos[13682]=-53;
cos[13683]=-53;
cos[13684]=-53;
cos[13685]=-53;
cos[13686]=-53;
cos[13687]=-53;
cos[13688]=-53;
cos[13689]=-53;
cos[13690]=-53;
cos[13691]=-53;
cos[13692]=-53;
cos[13693]=-53;
cos[13694]=-53;
cos[13695]=-53;
cos[13696]=-53;
cos[13697]=-53;
cos[13698]=-53;
cos[13699]=-53;
cos[13700]=-53;
cos[13701]=-54;
cos[13702]=-54;
cos[13703]=-54;
cos[13704]=-54;
cos[13705]=-54;
cos[13706]=-54;
cos[13707]=-54;
cos[13708]=-54;
cos[13709]=-54;
cos[13710]=-54;
cos[13711]=-54;
cos[13712]=-54;
cos[13713]=-54;
cos[13714]=-54;
cos[13715]=-54;
cos[13716]=-54;
cos[13717]=-54;
cos[13718]=-54;
cos[13719]=-54;
cos[13720]=-54;
cos[13721]=-54;
cos[13722]=-54;
cos[13723]=-54;
cos[13724]=-54;
cos[13725]=-54;
cos[13726]=-54;
cos[13727]=-54;
cos[13728]=-54;
cos[13729]=-55;
cos[13730]=-55;
cos[13731]=-55;
cos[13732]=-55;
cos[13733]=-55;
cos[13734]=-55;
cos[13735]=-55;
cos[13736]=-55;
cos[13737]=-55;
cos[13738]=-55;
cos[13739]=-55;
cos[13740]=-55;
cos[13741]=-55;
cos[13742]=-55;
cos[13743]=-55;
cos[13744]=-55;
cos[13745]=-55;
cos[13746]=-55;
cos[13747]=-55;
cos[13748]=-55;
cos[13749]=-55;
cos[13750]=-55;
cos[13751]=-55;
cos[13752]=-55;
cos[13753]=-55;
cos[13754]=-55;
cos[13755]=-55;
cos[13756]=-55;
cos[13757]=-55;
cos[13758]=-56;
cos[13759]=-56;
cos[13760]=-56;
cos[13761]=-56;
cos[13762]=-56;
cos[13763]=-56;
cos[13764]=-56;
cos[13765]=-56;
cos[13766]=-56;
cos[13767]=-56;
cos[13768]=-56;
cos[13769]=-56;
cos[13770]=-56;
cos[13771]=-56;
cos[13772]=-56;
cos[13773]=-56;
cos[13774]=-56;
cos[13775]=-56;
cos[13776]=-56;
cos[13777]=-56;
cos[13778]=-56;
cos[13779]=-56;
cos[13780]=-56;
cos[13781]=-56;
cos[13782]=-56;
cos[13783]=-56;
cos[13784]=-56;
cos[13785]=-56;
cos[13786]=-56;
cos[13787]=-57;
cos[13788]=-57;
cos[13789]=-57;
cos[13790]=-57;
cos[13791]=-57;
cos[13792]=-57;
cos[13793]=-57;
cos[13794]=-57;
cos[13795]=-57;
cos[13796]=-57;
cos[13797]=-57;
cos[13798]=-57;
cos[13799]=-57;
cos[13800]=-57;
cos[13801]=-57;
cos[13802]=-57;
cos[13803]=-57;
cos[13804]=-57;
cos[13805]=-57;
cos[13806]=-57;
cos[13807]=-57;
cos[13808]=-57;
cos[13809]=-57;
cos[13810]=-57;
cos[13811]=-57;
cos[13812]=-57;
cos[13813]=-57;
cos[13814]=-57;
cos[13815]=-57;
cos[13816]=-57;
cos[13817]=-58;
cos[13818]=-58;
cos[13819]=-58;
cos[13820]=-58;
cos[13821]=-58;
cos[13822]=-58;
cos[13823]=-58;
cos[13824]=-58;
cos[13825]=-58;
cos[13826]=-58;
cos[13827]=-58;
cos[13828]=-58;
cos[13829]=-58;
cos[13830]=-58;
cos[13831]=-58;
cos[13832]=-58;
cos[13833]=-58;
cos[13834]=-58;
cos[13835]=-58;
cos[13836]=-58;
cos[13837]=-58;
cos[13838]=-58;
cos[13839]=-58;
cos[13840]=-58;
cos[13841]=-58;
cos[13842]=-58;
cos[13843]=-58;
cos[13844]=-58;
cos[13845]=-58;
cos[13846]=-58;
cos[13847]=-59;
cos[13848]=-59;
cos[13849]=-59;
cos[13850]=-59;
cos[13851]=-59;
cos[13852]=-59;
cos[13853]=-59;
cos[13854]=-59;
cos[13855]=-59;
cos[13856]=-59;
cos[13857]=-59;
cos[13858]=-59;
cos[13859]=-59;
cos[13860]=-59;
cos[13861]=-59;
cos[13862]=-59;
cos[13863]=-59;
cos[13864]=-59;
cos[13865]=-59;
cos[13866]=-59;
cos[13867]=-59;
cos[13868]=-59;
cos[13869]=-59;
cos[13870]=-59;
cos[13871]=-59;
cos[13872]=-59;
cos[13873]=-59;
cos[13874]=-59;
cos[13875]=-59;
cos[13876]=-59;
cos[13877]=-59;
cos[13878]=-60;
cos[13879]=-60;
cos[13880]=-60;
cos[13881]=-60;
cos[13882]=-60;
cos[13883]=-60;
cos[13884]=-60;
cos[13885]=-60;
cos[13886]=-60;
cos[13887]=-60;
cos[13888]=-60;
cos[13889]=-60;
cos[13890]=-60;
cos[13891]=-60;
cos[13892]=-60;
cos[13893]=-60;
cos[13894]=-60;
cos[13895]=-60;
cos[13896]=-60;
cos[13897]=-60;
cos[13898]=-60;
cos[13899]=-60;
cos[13900]=-60;
cos[13901]=-60;
cos[13902]=-60;
cos[13903]=-60;
cos[13904]=-60;
cos[13905]=-60;
cos[13906]=-60;
cos[13907]=-60;
cos[13908]=-60;
cos[13909]=-60;
cos[13910]=-61;
cos[13911]=-61;
cos[13912]=-61;
cos[13913]=-61;
cos[13914]=-61;
cos[13915]=-61;
cos[13916]=-61;
cos[13917]=-61;
cos[13918]=-61;
cos[13919]=-61;
cos[13920]=-61;
cos[13921]=-61;
cos[13922]=-61;
cos[13923]=-61;
cos[13924]=-61;
cos[13925]=-61;
cos[13926]=-61;
cos[13927]=-61;
cos[13928]=-61;
cos[13929]=-61;
cos[13930]=-61;
cos[13931]=-61;
cos[13932]=-61;
cos[13933]=-61;
cos[13934]=-61;
cos[13935]=-61;
cos[13936]=-61;
cos[13937]=-61;
cos[13938]=-61;
cos[13939]=-61;
cos[13940]=-61;
cos[13941]=-61;
cos[13942]=-61;
cos[13943]=-62;
cos[13944]=-62;
cos[13945]=-62;
cos[13946]=-62;
cos[13947]=-62;
cos[13948]=-62;
cos[13949]=-62;
cos[13950]=-62;
cos[13951]=-62;
cos[13952]=-62;
cos[13953]=-62;
cos[13954]=-62;
cos[13955]=-62;
cos[13956]=-62;
cos[13957]=-62;
cos[13958]=-62;
cos[13959]=-62;
cos[13960]=-62;
cos[13961]=-62;
cos[13962]=-62;
cos[13963]=-62;
cos[13964]=-62;
cos[13965]=-62;
cos[13966]=-62;
cos[13967]=-62;
cos[13968]=-62;
cos[13969]=-62;
cos[13970]=-62;
cos[13971]=-62;
cos[13972]=-62;
cos[13973]=-62;
cos[13974]=-62;
cos[13975]=-62;
cos[13976]=-63;
cos[13977]=-63;
cos[13978]=-63;
cos[13979]=-63;
cos[13980]=-63;
cos[13981]=-63;
cos[13982]=-63;
cos[13983]=-63;
cos[13984]=-63;
cos[13985]=-63;
cos[13986]=-63;
cos[13987]=-63;
cos[13988]=-63;
cos[13989]=-63;
cos[13990]=-63;
cos[13991]=-63;
cos[13992]=-63;
cos[13993]=-63;
cos[13994]=-63;
cos[13995]=-63;
cos[13996]=-63;
cos[13997]=-63;
cos[13998]=-63;
cos[13999]=-63;
cos[14000]=-63;
cos[14001]=-63;
cos[14002]=-63;
cos[14003]=-63;
cos[14004]=-63;
cos[14005]=-63;
cos[14006]=-63;
cos[14007]=-63;
cos[14008]=-63;
cos[14009]=-63;
cos[14010]=-63;
cos[14011]=-64;
cos[14012]=-64;
cos[14013]=-64;
cos[14014]=-64;
cos[14015]=-64;
cos[14016]=-64;
cos[14017]=-64;
cos[14018]=-64;
cos[14019]=-64;
cos[14020]=-64;
cos[14021]=-64;
cos[14022]=-64;
cos[14023]=-64;
cos[14024]=-64;
cos[14025]=-64;
cos[14026]=-64;
cos[14027]=-64;
cos[14028]=-64;
cos[14029]=-64;
cos[14030]=-64;
cos[14031]=-64;
cos[14032]=-64;
cos[14033]=-64;
cos[14034]=-64;
cos[14035]=-64;
cos[14036]=-64;
cos[14037]=-64;
cos[14038]=-64;
cos[14039]=-64;
cos[14040]=-64;
cos[14041]=-64;
cos[14042]=-64;
cos[14043]=-64;
cos[14044]=-64;
cos[14045]=-64;
cos[14046]=-65;
cos[14047]=-65;
cos[14048]=-65;
cos[14049]=-65;
cos[14050]=-65;
cos[14051]=-65;
cos[14052]=-65;
cos[14053]=-65;
cos[14054]=-65;
cos[14055]=-65;
cos[14056]=-65;
cos[14057]=-65;
cos[14058]=-65;
cos[14059]=-65;
cos[14060]=-65;
cos[14061]=-65;
cos[14062]=-65;
cos[14063]=-65;
cos[14064]=-65;
cos[14065]=-65;
cos[14066]=-65;
cos[14067]=-65;
cos[14068]=-65;
cos[14069]=-65;
cos[14070]=-65;
cos[14071]=-65;
cos[14072]=-65;
cos[14073]=-65;
cos[14074]=-65;
cos[14075]=-65;
cos[14076]=-65;
cos[14077]=-65;
cos[14078]=-65;
cos[14079]=-65;
cos[14080]=-65;
cos[14081]=-65;
cos[14082]=-65;
cos[14083]=-66;
cos[14084]=-66;
cos[14085]=-66;
cos[14086]=-66;
cos[14087]=-66;
cos[14088]=-66;
cos[14089]=-66;
cos[14090]=-66;
cos[14091]=-66;
cos[14092]=-66;
cos[14093]=-66;
cos[14094]=-66;
cos[14095]=-66;
cos[14096]=-66;
cos[14097]=-66;
cos[14098]=-66;
cos[14099]=-66;
cos[14100]=-66;
cos[14101]=-66;
cos[14102]=-66;
cos[14103]=-66;
cos[14104]=-66;
cos[14105]=-66;
cos[14106]=-66;
cos[14107]=-66;
cos[14108]=-66;
cos[14109]=-66;
cos[14110]=-66;
cos[14111]=-66;
cos[14112]=-66;
cos[14113]=-66;
cos[14114]=-66;
cos[14115]=-66;
cos[14116]=-66;
cos[14117]=-66;
cos[14118]=-66;
cos[14119]=-66;
cos[14120]=-66;
cos[14121]=-67;
cos[14122]=-67;
cos[14123]=-67;
cos[14124]=-67;
cos[14125]=-67;
cos[14126]=-67;
cos[14127]=-67;
cos[14128]=-67;
cos[14129]=-67;
cos[14130]=-67;
cos[14131]=-67;
cos[14132]=-67;
cos[14133]=-67;
cos[14134]=-67;
cos[14135]=-67;
cos[14136]=-67;
cos[14137]=-67;
cos[14138]=-67;
cos[14139]=-67;
cos[14140]=-67;
cos[14141]=-67;
cos[14142]=-67;
cos[14143]=-67;
cos[14144]=-67;
cos[14145]=-67;
cos[14146]=-67;
cos[14147]=-67;
cos[14148]=-67;
cos[14149]=-67;
cos[14150]=-67;
cos[14151]=-67;
cos[14152]=-67;
cos[14153]=-67;
cos[14154]=-67;
cos[14155]=-67;
cos[14156]=-67;
cos[14157]=-67;
cos[14158]=-67;
cos[14159]=-67;
cos[14160]=-67;
cos[14161]=-68;
cos[14162]=-68;
cos[14163]=-68;
cos[14164]=-68;
cos[14165]=-68;
cos[14166]=-68;
cos[14167]=-68;
cos[14168]=-68;
cos[14169]=-68;
cos[14170]=-68;
cos[14171]=-68;
cos[14172]=-68;
cos[14173]=-68;
cos[14174]=-68;
cos[14175]=-68;
cos[14176]=-68;
cos[14177]=-68;
cos[14178]=-68;
cos[14179]=-68;
cos[14180]=-68;
cos[14181]=-68;
cos[14182]=-68;
cos[14183]=-68;
cos[14184]=-68;
cos[14185]=-68;
cos[14186]=-68;
cos[14187]=-68;
cos[14188]=-68;
cos[14189]=-68;
cos[14190]=-68;
cos[14191]=-68;
cos[14192]=-68;
cos[14193]=-68;
cos[14194]=-68;
cos[14195]=-68;
cos[14196]=-68;
cos[14197]=-68;
cos[14198]=-68;
cos[14199]=-68;
cos[14200]=-68;
cos[14201]=-68;
cos[14202]=-69;
cos[14203]=-69;
cos[14204]=-69;
cos[14205]=-69;
cos[14206]=-69;
cos[14207]=-69;
cos[14208]=-69;
cos[14209]=-69;
cos[14210]=-69;
cos[14211]=-69;
cos[14212]=-69;
cos[14213]=-69;
cos[14214]=-69;
cos[14215]=-69;
cos[14216]=-69;
cos[14217]=-69;
cos[14218]=-69;
cos[14219]=-69;
cos[14220]=-69;
cos[14221]=-69;
cos[14222]=-69;
cos[14223]=-69;
cos[14224]=-69;
cos[14225]=-69;
cos[14226]=-69;
cos[14227]=-69;
cos[14228]=-69;
cos[14229]=-69;
cos[14230]=-69;
cos[14231]=-69;
cos[14232]=-69;
cos[14233]=-69;
cos[14234]=-69;
cos[14235]=-69;
cos[14236]=-69;
cos[14237]=-69;
cos[14238]=-69;
cos[14239]=-69;
cos[14240]=-69;
cos[14241]=-69;
cos[14242]=-69;
cos[14243]=-69;
cos[14244]=-69;
cos[14245]=-69;
cos[14246]=-70;
cos[14247]=-70;
cos[14248]=-70;
cos[14249]=-70;
cos[14250]=-70;
cos[14251]=-70;
cos[14252]=-70;
cos[14253]=-70;
cos[14254]=-70;
cos[14255]=-70;
cos[14256]=-70;
cos[14257]=-70;
cos[14258]=-70;
cos[14259]=-70;
cos[14260]=-70;
cos[14261]=-70;
cos[14262]=-70;
cos[14263]=-70;
cos[14264]=-70;
cos[14265]=-70;
cos[14266]=-70;
cos[14267]=-70;
cos[14268]=-70;
cos[14269]=-70;
cos[14270]=-70;
cos[14271]=-70;
cos[14272]=-70;
cos[14273]=-70;
cos[14274]=-70;
cos[14275]=-70;
cos[14276]=-70;
cos[14277]=-70;
cos[14278]=-70;
cos[14279]=-70;
cos[14280]=-70;
cos[14281]=-70;
cos[14282]=-70;
cos[14283]=-70;
cos[14284]=-70;
cos[14285]=-70;
cos[14286]=-70;
cos[14287]=-70;
cos[14288]=-70;
cos[14289]=-70;
cos[14290]=-70;
cos[14291]=-71;
cos[14292]=-71;
cos[14293]=-71;
cos[14294]=-71;
cos[14295]=-71;
cos[14296]=-71;
cos[14297]=-71;
cos[14298]=-71;
cos[14299]=-71;
cos[14300]=-71;
cos[14301]=-71;
cos[14302]=-71;
cos[14303]=-71;
cos[14304]=-71;
cos[14305]=-71;
cos[14306]=-71;
cos[14307]=-71;
cos[14308]=-71;
cos[14309]=-71;
cos[14310]=-71;
cos[14311]=-71;
cos[14312]=-71;
cos[14313]=-71;
cos[14314]=-71;
cos[14315]=-71;
cos[14316]=-71;
cos[14317]=-71;
cos[14318]=-71;
cos[14319]=-71;
cos[14320]=-71;
cos[14321]=-71;
cos[14322]=-71;
cos[14323]=-71;
cos[14324]=-71;
cos[14325]=-71;
cos[14326]=-71;
cos[14327]=-71;
cos[14328]=-71;
cos[14329]=-71;
cos[14330]=-71;
cos[14331]=-71;
cos[14332]=-71;
cos[14333]=-71;
cos[14334]=-71;
cos[14335]=-71;
cos[14336]=-71;
cos[14337]=-71;
cos[14338]=-71;
cos[14339]=-71;
cos[14340]=-72;
cos[14341]=-72;
cos[14342]=-72;
cos[14343]=-72;
cos[14344]=-72;
cos[14345]=-72;
cos[14346]=-72;
cos[14347]=-72;
cos[14348]=-72;
cos[14349]=-72;
cos[14350]=-72;
cos[14351]=-72;
cos[14352]=-72;
cos[14353]=-72;
cos[14354]=-72;
cos[14355]=-72;
cos[14356]=-72;
cos[14357]=-72;
cos[14358]=-72;
cos[14359]=-72;
cos[14360]=-72;
cos[14361]=-72;
cos[14362]=-72;
cos[14363]=-72;
cos[14364]=-72;
cos[14365]=-72;
cos[14366]=-72;
cos[14367]=-72;
cos[14368]=-72;
cos[14369]=-72;
cos[14370]=-72;
cos[14371]=-72;
cos[14372]=-72;
cos[14373]=-72;
cos[14374]=-72;
cos[14375]=-72;
cos[14376]=-72;
cos[14377]=-72;
cos[14378]=-72;
cos[14379]=-72;
cos[14380]=-72;
cos[14381]=-72;
cos[14382]=-72;
cos[14383]=-72;
cos[14384]=-72;
cos[14385]=-72;
cos[14386]=-72;
cos[14387]=-72;
cos[14388]=-72;
cos[14389]=-72;
cos[14390]=-72;
cos[14391]=-72;
cos[14392]=-72;
cos[14393]=-73;
cos[14394]=-73;
cos[14395]=-73;
cos[14396]=-73;
cos[14397]=-73;
cos[14398]=-73;
cos[14399]=-73;
cos[14400]=-73;
cos[14401]=-73;
cos[14402]=-73;
cos[14403]=-73;
cos[14404]=-73;
cos[14405]=-73;
cos[14406]=-73;
cos[14407]=-73;
cos[14408]=-73;
cos[14409]=-73;
cos[14410]=-73;
cos[14411]=-73;
cos[14412]=-73;
cos[14413]=-73;
cos[14414]=-73;
cos[14415]=-73;
cos[14416]=-73;
cos[14417]=-73;
cos[14418]=-73;
cos[14419]=-73;
cos[14420]=-73;
cos[14421]=-73;
cos[14422]=-73;
cos[14423]=-73;
cos[14424]=-73;
cos[14425]=-73;
cos[14426]=-73;
cos[14427]=-73;
cos[14428]=-73;
cos[14429]=-73;
cos[14430]=-73;
cos[14431]=-73;
cos[14432]=-73;
cos[14433]=-73;
cos[14434]=-73;
cos[14435]=-73;
cos[14436]=-73;
cos[14437]=-73;
cos[14438]=-73;
cos[14439]=-73;
cos[14440]=-73;
cos[14441]=-73;
cos[14442]=-73;
cos[14443]=-73;
cos[14444]=-73;
cos[14445]=-73;
cos[14446]=-73;
cos[14447]=-73;
cos[14448]=-73;
cos[14449]=-73;
cos[14450]=-74;
cos[14451]=-74;
cos[14452]=-74;
cos[14453]=-74;
cos[14454]=-74;
cos[14455]=-74;
cos[14456]=-74;
cos[14457]=-74;
cos[14458]=-74;
cos[14459]=-74;
cos[14460]=-74;
cos[14461]=-74;
cos[14462]=-74;
cos[14463]=-74;
cos[14464]=-74;
cos[14465]=-74;
cos[14466]=-74;
cos[14467]=-74;
cos[14468]=-74;
cos[14469]=-74;
cos[14470]=-74;
cos[14471]=-74;
cos[14472]=-74;
cos[14473]=-74;
cos[14474]=-74;
cos[14475]=-74;
cos[14476]=-74;
cos[14477]=-74;
cos[14478]=-74;
cos[14479]=-74;
cos[14480]=-74;
cos[14481]=-74;
cos[14482]=-74;
cos[14483]=-74;
cos[14484]=-74;
cos[14485]=-74;
cos[14486]=-74;
cos[14487]=-74;
cos[14488]=-74;
cos[14489]=-74;
cos[14490]=-74;
cos[14491]=-74;
cos[14492]=-74;
cos[14493]=-74;
cos[14494]=-74;
cos[14495]=-74;
cos[14496]=-74;
cos[14497]=-74;
cos[14498]=-74;
cos[14499]=-74;
cos[14500]=-74;
cos[14501]=-74;
cos[14502]=-74;
cos[14503]=-74;
cos[14504]=-74;
cos[14505]=-74;
cos[14506]=-74;
cos[14507]=-74;
cos[14508]=-74;
cos[14509]=-74;
cos[14510]=-74;
cos[14511]=-74;
cos[14512]=-74;
cos[14513]=-74;
cos[14514]=-75;
cos[14515]=-75;
cos[14516]=-75;
cos[14517]=-75;
cos[14518]=-75;
cos[14519]=-75;
cos[14520]=-75;
cos[14521]=-75;
cos[14522]=-75;
cos[14523]=-75;
cos[14524]=-75;
cos[14525]=-75;
cos[14526]=-75;
cos[14527]=-75;
cos[14528]=-75;
cos[14529]=-75;
cos[14530]=-75;
cos[14531]=-75;
cos[14532]=-75;
cos[14533]=-75;
cos[14534]=-75;
cos[14535]=-75;
cos[14536]=-75;
cos[14537]=-75;
cos[14538]=-75;
cos[14539]=-75;
cos[14540]=-75;
cos[14541]=-75;
cos[14542]=-75;
cos[14543]=-75;
cos[14544]=-75;
cos[14545]=-75;
cos[14546]=-75;
cos[14547]=-75;
cos[14548]=-75;
cos[14549]=-75;
cos[14550]=-75;
cos[14551]=-75;
cos[14552]=-75;
cos[14553]=-75;
cos[14554]=-75;
cos[14555]=-75;
cos[14556]=-75;
cos[14557]=-75;
cos[14558]=-75;
cos[14559]=-75;
cos[14560]=-75;
cos[14561]=-75;
cos[14562]=-75;
cos[14563]=-75;
cos[14564]=-75;
cos[14565]=-75;
cos[14566]=-75;
cos[14567]=-75;
cos[14568]=-75;
cos[14569]=-75;
cos[14570]=-75;
cos[14571]=-75;
cos[14572]=-75;
cos[14573]=-75;
cos[14574]=-75;
cos[14575]=-75;
cos[14576]=-75;
cos[14577]=-75;
cos[14578]=-75;
cos[14579]=-75;
cos[14580]=-75;
cos[14581]=-75;
cos[14582]=-75;
cos[14583]=-75;
cos[14584]=-75;
cos[14585]=-75;
cos[14586]=-75;
cos[14587]=-76;
cos[14588]=-76;
cos[14589]=-76;
cos[14590]=-76;
cos[14591]=-76;
cos[14592]=-76;
cos[14593]=-76;
cos[14594]=-76;
cos[14595]=-76;
cos[14596]=-76;
cos[14597]=-76;
cos[14598]=-76;
cos[14599]=-76;
cos[14600]=-76;
cos[14601]=-76;
cos[14602]=-76;
cos[14603]=-76;
cos[14604]=-76;
cos[14605]=-76;
cos[14606]=-76;
cos[14607]=-76;
cos[14608]=-76;
cos[14609]=-76;
cos[14610]=-76;
cos[14611]=-76;
cos[14612]=-76;
cos[14613]=-76;
cos[14614]=-76;
cos[14615]=-76;
cos[14616]=-76;
cos[14617]=-76;
cos[14618]=-76;
cos[14619]=-76;
cos[14620]=-76;
cos[14621]=-76;
cos[14622]=-76;
cos[14623]=-76;
cos[14624]=-76;
cos[14625]=-76;
cos[14626]=-76;
cos[14627]=-76;
cos[14628]=-76;
cos[14629]=-76;
cos[14630]=-76;
cos[14631]=-76;
cos[14632]=-76;
cos[14633]=-76;
cos[14634]=-76;
cos[14635]=-76;
cos[14636]=-76;
cos[14637]=-76;
cos[14638]=-76;
cos[14639]=-76;
cos[14640]=-76;
cos[14641]=-76;
cos[14642]=-76;
cos[14643]=-76;
cos[14644]=-76;
cos[14645]=-76;
cos[14646]=-76;
cos[14647]=-76;
cos[14648]=-76;
cos[14649]=-76;
cos[14650]=-76;
cos[14651]=-76;
cos[14652]=-76;
cos[14653]=-76;
cos[14654]=-76;
cos[14655]=-76;
cos[14656]=-76;
cos[14657]=-76;
cos[14658]=-76;
cos[14659]=-76;
cos[14660]=-76;
cos[14661]=-76;
cos[14662]=-76;
cos[14663]=-76;
cos[14664]=-76;
cos[14665]=-76;
cos[14666]=-76;
cos[14667]=-76;
cos[14668]=-76;
cos[14669]=-76;
cos[14670]=-76;
cos[14671]=-76;
cos[14672]=-76;
cos[14673]=-76;
cos[14674]=-76;
cos[14675]=-77;
cos[14676]=-77;
cos[14677]=-77;
cos[14678]=-77;
cos[14679]=-77;
cos[14680]=-77;
cos[14681]=-77;
cos[14682]=-77;
cos[14683]=-77;
cos[14684]=-77;
cos[14685]=-77;
cos[14686]=-77;
cos[14687]=-77;
cos[14688]=-77;
cos[14689]=-77;
cos[14690]=-77;
cos[14691]=-77;
cos[14692]=-77;
cos[14693]=-77;
cos[14694]=-77;
cos[14695]=-77;
cos[14696]=-77;
cos[14697]=-77;
cos[14698]=-77;
cos[14699]=-77;
cos[14700]=-77;
cos[14701]=-77;
cos[14702]=-77;
cos[14703]=-77;
cos[14704]=-77;
cos[14705]=-77;
cos[14706]=-77;
cos[14707]=-77;
cos[14708]=-77;
cos[14709]=-77;
cos[14710]=-77;
cos[14711]=-77;
cos[14712]=-77;
cos[14713]=-77;
cos[14714]=-77;
cos[14715]=-77;
cos[14716]=-77;
cos[14717]=-77;
cos[14718]=-77;
cos[14719]=-77;
cos[14720]=-77;
cos[14721]=-77;
cos[14722]=-77;
cos[14723]=-77;
cos[14724]=-77;
cos[14725]=-77;
cos[14726]=-77;
cos[14727]=-77;
cos[14728]=-77;
cos[14729]=-77;
cos[14730]=-77;
cos[14731]=-77;
cos[14732]=-77;
cos[14733]=-77;
cos[14734]=-77;
cos[14735]=-77;
cos[14736]=-77;
cos[14737]=-77;
cos[14738]=-77;
cos[14739]=-77;
cos[14740]=-77;
cos[14741]=-77;
cos[14742]=-77;
cos[14743]=-77;
cos[14744]=-77;
cos[14745]=-77;
cos[14746]=-77;
cos[14747]=-77;
cos[14748]=-77;
cos[14749]=-77;
cos[14750]=-77;
cos[14751]=-77;
cos[14752]=-77;
cos[14753]=-77;
cos[14754]=-77;
cos[14755]=-77;
cos[14756]=-77;
cos[14757]=-77;
cos[14758]=-77;
cos[14759]=-77;
cos[14760]=-77;
cos[14761]=-77;
cos[14762]=-77;
cos[14763]=-77;
cos[14764]=-77;
cos[14765]=-77;
cos[14766]=-77;
cos[14767]=-77;
cos[14768]=-77;
cos[14769]=-77;
cos[14770]=-77;
cos[14771]=-77;
cos[14772]=-77;
cos[14773]=-77;
cos[14774]=-77;
cos[14775]=-77;
cos[14776]=-77;
cos[14777]=-77;
cos[14778]=-77;
cos[14779]=-77;
cos[14780]=-77;
cos[14781]=-77;
cos[14782]=-77;
cos[14783]=-77;
cos[14784]=-77;
cos[14785]=-77;
cos[14786]=-77;
cos[14787]=-77;
cos[14788]=-77;
cos[14789]=-77;
cos[14790]=-77;
cos[14791]=-77;
cos[14792]=-77;
cos[14793]=-77;
cos[14794]=-77;
cos[14795]=-77;
cos[14796]=-77;
cos[14797]=-77;
cos[14798]=-77;
cos[14799]=-78;
cos[14800]=-78;
cos[14801]=-78;
cos[14802]=-78;
cos[14803]=-78;
cos[14804]=-78;
cos[14805]=-78;
cos[14806]=-78;
cos[14807]=-78;
cos[14808]=-78;
cos[14809]=-78;
cos[14810]=-78;
cos[14811]=-78;
cos[14812]=-78;
cos[14813]=-78;
cos[14814]=-78;
cos[14815]=-78;
cos[14816]=-78;
cos[14817]=-78;
cos[14818]=-78;
cos[14819]=-78;
cos[14820]=-78;
cos[14821]=-78;
cos[14822]=-78;
cos[14823]=-78;
cos[14824]=-78;
cos[14825]=-78;
cos[14826]=-78;
cos[14827]=-78;
cos[14828]=-78;
cos[14829]=-78;
cos[14830]=-78;
cos[14831]=-78;
cos[14832]=-78;
cos[14833]=-78;
cos[14834]=-78;
cos[14835]=-78;
cos[14836]=-78;
cos[14837]=-78;
cos[14838]=-78;
cos[14839]=-78;
cos[14840]=-78;
cos[14841]=-78;
cos[14842]=-78;
cos[14843]=-78;
cos[14844]=-78;
cos[14845]=-78;
cos[14846]=-78;
cos[14847]=-78;
cos[14848]=-78;
cos[14849]=-78;
cos[14850]=-78;
cos[14851]=-78;
cos[14852]=-78;
cos[14853]=-78;
cos[14854]=-78;
cos[14855]=-78;
cos[14856]=-78;
cos[14857]=-78;
cos[14858]=-78;
cos[14859]=-78;
cos[14860]=-78;
cos[14861]=-78;
cos[14862]=-78;
cos[14863]=-78;
cos[14864]=-78;
cos[14865]=-78;
cos[14866]=-78;
cos[14867]=-78;
cos[14868]=-78;
cos[14869]=-78;
cos[14870]=-78;
cos[14871]=-78;
cos[14872]=-78;
cos[14873]=-78;
cos[14874]=-78;
cos[14875]=-78;
cos[14876]=-78;
cos[14877]=-78;
cos[14878]=-78;
cos[14879]=-78;
cos[14880]=-78;
cos[14881]=-78;
cos[14882]=-78;
cos[14883]=-78;
cos[14884]=-78;
cos[14885]=-78;
cos[14886]=-78;
cos[14887]=-78;
cos[14888]=-78;
cos[14889]=-78;
cos[14890]=-78;
cos[14891]=-78;
cos[14892]=-78;
cos[14893]=-78;
cos[14894]=-78;
cos[14895]=-78;
cos[14896]=-78;
cos[14897]=-78;
cos[14898]=-78;
cos[14899]=-78;
cos[14900]=-78;
cos[14901]=-78;
cos[14902]=-78;
cos[14903]=-78;
cos[14904]=-78;
cos[14905]=-78;
cos[14906]=-78;
cos[14907]=-78;
cos[14908]=-78;
cos[14909]=-78;
cos[14910]=-78;
cos[14911]=-78;
cos[14912]=-78;
cos[14913]=-78;
cos[14914]=-78;
cos[14915]=-78;
cos[14916]=-78;
cos[14917]=-78;
cos[14918]=-78;
cos[14919]=-78;
cos[14920]=-78;
cos[14921]=-78;
cos[14922]=-78;
cos[14923]=-78;
cos[14924]=-78;
cos[14925]=-78;
cos[14926]=-78;
cos[14927]=-78;
cos[14928]=-78;
cos[14929]=-78;
cos[14930]=-78;
cos[14931]=-78;
cos[14932]=-78;
cos[14933]=-78;
cos[14934]=-78;
cos[14935]=-78;
cos[14936]=-78;
cos[14937]=-78;
cos[14938]=-78;
cos[14939]=-78;
cos[14940]=-78;
cos[14941]=-78;
cos[14942]=-78;
cos[14943]=-78;
cos[14944]=-78;
cos[14945]=-78;
cos[14946]=-78;
cos[14947]=-78;
cos[14948]=-78;
cos[14949]=-78;
cos[14950]=-78;
cos[14951]=-78;
cos[14952]=-78;
cos[14953]=-78;
cos[14954]=-78;
cos[14955]=-78;
cos[14956]=-78;
cos[14957]=-78;
cos[14958]=-78;
cos[14959]=-78;
cos[14960]=-78;
cos[14961]=-78;
cos[14962]=-78;
cos[14963]=-78;
cos[14964]=-78;
cos[14965]=-78;
cos[14966]=-78;
cos[14967]=-78;
cos[14968]=-78;
cos[14969]=-78;
cos[14970]=-78;
cos[14971]=-78;
cos[14972]=-78;
cos[14973]=-78;
cos[14974]=-78;
cos[14975]=-78;
cos[14976]=-78;
cos[14977]=-78;
cos[14978]=-78;
cos[14979]=-78;
cos[14980]=-78;
cos[14981]=-78;
cos[14982]=-78;
cos[14983]=-78;
cos[14984]=-78;
cos[14985]=-78;
cos[14986]=-78;
cos[14987]=-78;
cos[14988]=-78;
cos[14989]=-78;
cos[14990]=-78;
cos[14991]=-78;
cos[14992]=-78;
cos[14993]=-78;
cos[14994]=-78;
cos[14995]=-78;
cos[14996]=-78;
cos[14997]=-78;
cos[14998]=-78;
cos[14999]=-78;
cos[15000]=-78;
cos[15001]=-78;
cos[15002]=-78;
cos[15003]=-78;
cos[15004]=-78;
cos[15005]=-78;
cos[15006]=-78;
cos[15007]=-78;
cos[15008]=-78;
cos[15009]=-78;
cos[15010]=-78;
cos[15011]=-78;
cos[15012]=-78;
cos[15013]=-78;
cos[15014]=-78;
cos[15015]=-78;
cos[15016]=-78;
cos[15017]=-78;
cos[15018]=-78;
cos[15019]=-78;
cos[15020]=-78;
cos[15021]=-78;
cos[15022]=-78;
cos[15023]=-78;
cos[15024]=-78;
cos[15025]=-78;
cos[15026]=-78;
cos[15027]=-78;
cos[15028]=-78;
cos[15029]=-78;
cos[15030]=-78;
cos[15031]=-78;
cos[15032]=-78;
cos[15033]=-78;
cos[15034]=-78;
cos[15035]=-78;
cos[15036]=-78;
cos[15037]=-78;
cos[15038]=-78;
cos[15039]=-78;
cos[15040]=-78;
cos[15041]=-78;
cos[15042]=-78;
cos[15043]=-78;
cos[15044]=-78;
cos[15045]=-78;
cos[15046]=-78;
cos[15047]=-78;
cos[15048]=-78;
cos[15049]=-78;
cos[15050]=-78;
cos[15051]=-78;
cos[15052]=-78;
cos[15053]=-78;
cos[15054]=-78;
cos[15055]=-78;
cos[15056]=-78;
cos[15057]=-78;
cos[15058]=-78;
cos[15059]=-78;
cos[15060]=-78;
cos[15061]=-78;
cos[15062]=-78;
cos[15063]=-78;
cos[15064]=-78;
cos[15065]=-78;
cos[15066]=-78;
cos[15067]=-78;
cos[15068]=-78;
cos[15069]=-78;
cos[15070]=-78;
cos[15071]=-78;
cos[15072]=-78;
cos[15073]=-78;
cos[15074]=-78;
cos[15075]=-78;
cos[15076]=-78;
cos[15077]=-78;
cos[15078]=-78;
cos[15079]=-78;
cos[15080]=-78;
cos[15081]=-78;
cos[15082]=-78;
cos[15083]=-78;
cos[15084]=-78;
cos[15085]=-78;
cos[15086]=-78;
cos[15087]=-78;
cos[15088]=-78;
cos[15089]=-78;
cos[15090]=-78;
cos[15091]=-78;
cos[15092]=-78;
cos[15093]=-78;
cos[15094]=-78;
cos[15095]=-78;
cos[15096]=-78;
cos[15097]=-78;
cos[15098]=-78;
cos[15099]=-78;
cos[15100]=-78;
cos[15101]=-78;
cos[15102]=-78;
cos[15103]=-78;
cos[15104]=-78;
cos[15105]=-78;
cos[15106]=-78;
cos[15107]=-78;
cos[15108]=-78;
cos[15109]=-78;
cos[15110]=-78;
cos[15111]=-78;
cos[15112]=-78;
cos[15113]=-78;
cos[15114]=-78;
cos[15115]=-78;
cos[15116]=-78;
cos[15117]=-78;
cos[15118]=-78;
cos[15119]=-78;
cos[15120]=-78;
cos[15121]=-78;
cos[15122]=-78;
cos[15123]=-78;
cos[15124]=-78;
cos[15125]=-78;
cos[15126]=-78;
cos[15127]=-78;
cos[15128]=-78;
cos[15129]=-78;
cos[15130]=-78;
cos[15131]=-78;
cos[15132]=-78;
cos[15133]=-78;
cos[15134]=-78;
cos[15135]=-78;
cos[15136]=-78;
cos[15137]=-78;
cos[15138]=-78;
cos[15139]=-78;
cos[15140]=-78;
cos[15141]=-78;
cos[15142]=-78;
cos[15143]=-78;
cos[15144]=-78;
cos[15145]=-78;
cos[15146]=-78;
cos[15147]=-78;
cos[15148]=-78;
cos[15149]=-78;
cos[15150]=-78;
cos[15151]=-78;
cos[15152]=-78;
cos[15153]=-78;
cos[15154]=-78;
cos[15155]=-78;
cos[15156]=-78;
cos[15157]=-78;
cos[15158]=-78;
cos[15159]=-78;
cos[15160]=-78;
cos[15161]=-78;
cos[15162]=-78;
cos[15163]=-78;
cos[15164]=-78;
cos[15165]=-78;
cos[15166]=-78;
cos[15167]=-78;
cos[15168]=-78;
cos[15169]=-78;
cos[15170]=-78;
cos[15171]=-78;
cos[15172]=-78;
cos[15173]=-78;
cos[15174]=-78;
cos[15175]=-78;
cos[15176]=-78;
cos[15177]=-78;
cos[15178]=-78;
cos[15179]=-78;
cos[15180]=-78;
cos[15181]=-78;
cos[15182]=-78;
cos[15183]=-78;
cos[15184]=-78;
cos[15185]=-78;
cos[15186]=-78;
cos[15187]=-78;
cos[15188]=-78;
cos[15189]=-78;
cos[15190]=-78;
cos[15191]=-78;
cos[15192]=-78;
cos[15193]=-78;
cos[15194]=-78;
cos[15195]=-78;
cos[15196]=-78;
cos[15197]=-78;
cos[15198]=-78;
cos[15199]=-78;
cos[15200]=-78;
cos[15201]=-78;
cos[15202]=-77;
cos[15203]=-77;
cos[15204]=-77;
cos[15205]=-77;
cos[15206]=-77;
cos[15207]=-77;
cos[15208]=-77;
cos[15209]=-77;
cos[15210]=-77;
cos[15211]=-77;
cos[15212]=-77;
cos[15213]=-77;
cos[15214]=-77;
cos[15215]=-77;
cos[15216]=-77;
cos[15217]=-77;
cos[15218]=-77;
cos[15219]=-77;
cos[15220]=-77;
cos[15221]=-77;
cos[15222]=-77;
cos[15223]=-77;
cos[15224]=-77;
cos[15225]=-77;
cos[15226]=-77;
cos[15227]=-77;
cos[15228]=-77;
cos[15229]=-77;
cos[15230]=-77;
cos[15231]=-77;
cos[15232]=-77;
cos[15233]=-77;
cos[15234]=-77;
cos[15235]=-77;
cos[15236]=-77;
cos[15237]=-77;
cos[15238]=-77;
cos[15239]=-77;
cos[15240]=-77;
cos[15241]=-77;
cos[15242]=-77;
cos[15243]=-77;
cos[15244]=-77;
cos[15245]=-77;
cos[15246]=-77;
cos[15247]=-77;
cos[15248]=-77;
cos[15249]=-77;
cos[15250]=-77;
cos[15251]=-77;
cos[15252]=-77;
cos[15253]=-77;
cos[15254]=-77;
cos[15255]=-77;
cos[15256]=-77;
cos[15257]=-77;
cos[15258]=-77;
cos[15259]=-77;
cos[15260]=-77;
cos[15261]=-77;
cos[15262]=-77;
cos[15263]=-77;
cos[15264]=-77;
cos[15265]=-77;
cos[15266]=-77;
cos[15267]=-77;
cos[15268]=-77;
cos[15269]=-77;
cos[15270]=-77;
cos[15271]=-77;
cos[15272]=-77;
cos[15273]=-77;
cos[15274]=-77;
cos[15275]=-77;
cos[15276]=-77;
cos[15277]=-77;
cos[15278]=-77;
cos[15279]=-77;
cos[15280]=-77;
cos[15281]=-77;
cos[15282]=-77;
cos[15283]=-77;
cos[15284]=-77;
cos[15285]=-77;
cos[15286]=-77;
cos[15287]=-77;
cos[15288]=-77;
cos[15289]=-77;
cos[15290]=-77;
cos[15291]=-77;
cos[15292]=-77;
cos[15293]=-77;
cos[15294]=-77;
cos[15295]=-77;
cos[15296]=-77;
cos[15297]=-77;
cos[15298]=-77;
cos[15299]=-77;
cos[15300]=-77;
cos[15301]=-77;
cos[15302]=-77;
cos[15303]=-77;
cos[15304]=-77;
cos[15305]=-77;
cos[15306]=-77;
cos[15307]=-77;
cos[15308]=-77;
cos[15309]=-77;
cos[15310]=-77;
cos[15311]=-77;
cos[15312]=-77;
cos[15313]=-77;
cos[15314]=-77;
cos[15315]=-77;
cos[15316]=-77;
cos[15317]=-77;
cos[15318]=-77;
cos[15319]=-77;
cos[15320]=-77;
cos[15321]=-77;
cos[15322]=-77;
cos[15323]=-77;
cos[15324]=-77;
cos[15325]=-77;
cos[15326]=-76;
cos[15327]=-76;
cos[15328]=-76;
cos[15329]=-76;
cos[15330]=-76;
cos[15331]=-76;
cos[15332]=-76;
cos[15333]=-76;
cos[15334]=-76;
cos[15335]=-76;
cos[15336]=-76;
cos[15337]=-76;
cos[15338]=-76;
cos[15339]=-76;
cos[15340]=-76;
cos[15341]=-76;
cos[15342]=-76;
cos[15343]=-76;
cos[15344]=-76;
cos[15345]=-76;
cos[15346]=-76;
cos[15347]=-76;
cos[15348]=-76;
cos[15349]=-76;
cos[15350]=-76;
cos[15351]=-76;
cos[15352]=-76;
cos[15353]=-76;
cos[15354]=-76;
cos[15355]=-76;
cos[15356]=-76;
cos[15357]=-76;
cos[15358]=-76;
cos[15359]=-76;
cos[15360]=-76;
cos[15361]=-76;
cos[15362]=-76;
cos[15363]=-76;
cos[15364]=-76;
cos[15365]=-76;
cos[15366]=-76;
cos[15367]=-76;
cos[15368]=-76;
cos[15369]=-76;
cos[15370]=-76;
cos[15371]=-76;
cos[15372]=-76;
cos[15373]=-76;
cos[15374]=-76;
cos[15375]=-76;
cos[15376]=-76;
cos[15377]=-76;
cos[15378]=-76;
cos[15379]=-76;
cos[15380]=-76;
cos[15381]=-76;
cos[15382]=-76;
cos[15383]=-76;
cos[15384]=-76;
cos[15385]=-76;
cos[15386]=-76;
cos[15387]=-76;
cos[15388]=-76;
cos[15389]=-76;
cos[15390]=-76;
cos[15391]=-76;
cos[15392]=-76;
cos[15393]=-76;
cos[15394]=-76;
cos[15395]=-76;
cos[15396]=-76;
cos[15397]=-76;
cos[15398]=-76;
cos[15399]=-76;
cos[15400]=-76;
cos[15401]=-76;
cos[15402]=-76;
cos[15403]=-76;
cos[15404]=-76;
cos[15405]=-76;
cos[15406]=-76;
cos[15407]=-76;
cos[15408]=-76;
cos[15409]=-76;
cos[15410]=-76;
cos[15411]=-76;
cos[15412]=-76;
cos[15413]=-76;
cos[15414]=-75;
cos[15415]=-75;
cos[15416]=-75;
cos[15417]=-75;
cos[15418]=-75;
cos[15419]=-75;
cos[15420]=-75;
cos[15421]=-75;
cos[15422]=-75;
cos[15423]=-75;
cos[15424]=-75;
cos[15425]=-75;
cos[15426]=-75;
cos[15427]=-75;
cos[15428]=-75;
cos[15429]=-75;
cos[15430]=-75;
cos[15431]=-75;
cos[15432]=-75;
cos[15433]=-75;
cos[15434]=-75;
cos[15435]=-75;
cos[15436]=-75;
cos[15437]=-75;
cos[15438]=-75;
cos[15439]=-75;
cos[15440]=-75;
cos[15441]=-75;
cos[15442]=-75;
cos[15443]=-75;
cos[15444]=-75;
cos[15445]=-75;
cos[15446]=-75;
cos[15447]=-75;
cos[15448]=-75;
cos[15449]=-75;
cos[15450]=-75;
cos[15451]=-75;
cos[15452]=-75;
cos[15453]=-75;
cos[15454]=-75;
cos[15455]=-75;
cos[15456]=-75;
cos[15457]=-75;
cos[15458]=-75;
cos[15459]=-75;
cos[15460]=-75;
cos[15461]=-75;
cos[15462]=-75;
cos[15463]=-75;
cos[15464]=-75;
cos[15465]=-75;
cos[15466]=-75;
cos[15467]=-75;
cos[15468]=-75;
cos[15469]=-75;
cos[15470]=-75;
cos[15471]=-75;
cos[15472]=-75;
cos[15473]=-75;
cos[15474]=-75;
cos[15475]=-75;
cos[15476]=-75;
cos[15477]=-75;
cos[15478]=-75;
cos[15479]=-75;
cos[15480]=-75;
cos[15481]=-75;
cos[15482]=-75;
cos[15483]=-75;
cos[15484]=-75;
cos[15485]=-75;
cos[15486]=-75;
cos[15487]=-74;
cos[15488]=-74;
cos[15489]=-74;
cos[15490]=-74;
cos[15491]=-74;
cos[15492]=-74;
cos[15493]=-74;
cos[15494]=-74;
cos[15495]=-74;
cos[15496]=-74;
cos[15497]=-74;
cos[15498]=-74;
cos[15499]=-74;
cos[15500]=-74;
cos[15501]=-74;
cos[15502]=-74;
cos[15503]=-74;
cos[15504]=-74;
cos[15505]=-74;
cos[15506]=-74;
cos[15507]=-74;
cos[15508]=-74;
cos[15509]=-74;
cos[15510]=-74;
cos[15511]=-74;
cos[15512]=-74;
cos[15513]=-74;
cos[15514]=-74;
cos[15515]=-74;
cos[15516]=-74;
cos[15517]=-74;
cos[15518]=-74;
cos[15519]=-74;
cos[15520]=-74;
cos[15521]=-74;
cos[15522]=-74;
cos[15523]=-74;
cos[15524]=-74;
cos[15525]=-74;
cos[15526]=-74;
cos[15527]=-74;
cos[15528]=-74;
cos[15529]=-74;
cos[15530]=-74;
cos[15531]=-74;
cos[15532]=-74;
cos[15533]=-74;
cos[15534]=-74;
cos[15535]=-74;
cos[15536]=-74;
cos[15537]=-74;
cos[15538]=-74;
cos[15539]=-74;
cos[15540]=-74;
cos[15541]=-74;
cos[15542]=-74;
cos[15543]=-74;
cos[15544]=-74;
cos[15545]=-74;
cos[15546]=-74;
cos[15547]=-74;
cos[15548]=-74;
cos[15549]=-74;
cos[15550]=-74;
cos[15551]=-73;
cos[15552]=-73;
cos[15553]=-73;
cos[15554]=-73;
cos[15555]=-73;
cos[15556]=-73;
cos[15557]=-73;
cos[15558]=-73;
cos[15559]=-73;
cos[15560]=-73;
cos[15561]=-73;
cos[15562]=-73;
cos[15563]=-73;
cos[15564]=-73;
cos[15565]=-73;
cos[15566]=-73;
cos[15567]=-73;
cos[15568]=-73;
cos[15569]=-73;
cos[15570]=-73;
cos[15571]=-73;
cos[15572]=-73;
cos[15573]=-73;
cos[15574]=-73;
cos[15575]=-73;
cos[15576]=-73;
cos[15577]=-73;
cos[15578]=-73;
cos[15579]=-73;
cos[15580]=-73;
cos[15581]=-73;
cos[15582]=-73;
cos[15583]=-73;
cos[15584]=-73;
cos[15585]=-73;
cos[15586]=-73;
cos[15587]=-73;
cos[15588]=-73;
cos[15589]=-73;
cos[15590]=-73;
cos[15591]=-73;
cos[15592]=-73;
cos[15593]=-73;
cos[15594]=-73;
cos[15595]=-73;
cos[15596]=-73;
cos[15597]=-73;
cos[15598]=-73;
cos[15599]=-73;
cos[15600]=-73;
cos[15601]=-73;
cos[15602]=-73;
cos[15603]=-73;
cos[15604]=-73;
cos[15605]=-73;
cos[15606]=-73;
cos[15607]=-73;
cos[15608]=-72;
cos[15609]=-72;
cos[15610]=-72;
cos[15611]=-72;
cos[15612]=-72;
cos[15613]=-72;
cos[15614]=-72;
cos[15615]=-72;
cos[15616]=-72;
cos[15617]=-72;
cos[15618]=-72;
cos[15619]=-72;
cos[15620]=-72;
cos[15621]=-72;
cos[15622]=-72;
cos[15623]=-72;
cos[15624]=-72;
cos[15625]=-72;
cos[15626]=-72;
cos[15627]=-72;
cos[15628]=-72;
cos[15629]=-72;
cos[15630]=-72;
cos[15631]=-72;
cos[15632]=-72;
cos[15633]=-72;
cos[15634]=-72;
cos[15635]=-72;
cos[15636]=-72;
cos[15637]=-72;
cos[15638]=-72;
cos[15639]=-72;
cos[15640]=-72;
cos[15641]=-72;
cos[15642]=-72;
cos[15643]=-72;
cos[15644]=-72;
cos[15645]=-72;
cos[15646]=-72;
cos[15647]=-72;
cos[15648]=-72;
cos[15649]=-72;
cos[15650]=-72;
cos[15651]=-72;
cos[15652]=-72;
cos[15653]=-72;
cos[15654]=-72;
cos[15655]=-72;
cos[15656]=-72;
cos[15657]=-72;
cos[15658]=-72;
cos[15659]=-72;
cos[15660]=-72;
cos[15661]=-71;
cos[15662]=-71;
cos[15663]=-71;
cos[15664]=-71;
cos[15665]=-71;
cos[15666]=-71;
cos[15667]=-71;
cos[15668]=-71;
cos[15669]=-71;
cos[15670]=-71;
cos[15671]=-71;
cos[15672]=-71;
cos[15673]=-71;
cos[15674]=-71;
cos[15675]=-71;
cos[15676]=-71;
cos[15677]=-71;
cos[15678]=-71;
cos[15679]=-71;
cos[15680]=-71;
cos[15681]=-71;
cos[15682]=-71;
cos[15683]=-71;
cos[15684]=-71;
cos[15685]=-71;
cos[15686]=-71;
cos[15687]=-71;
cos[15688]=-71;
cos[15689]=-71;
cos[15690]=-71;
cos[15691]=-71;
cos[15692]=-71;
cos[15693]=-71;
cos[15694]=-71;
cos[15695]=-71;
cos[15696]=-71;
cos[15697]=-71;
cos[15698]=-71;
cos[15699]=-71;
cos[15700]=-71;
cos[15701]=-71;
cos[15702]=-71;
cos[15703]=-71;
cos[15704]=-71;
cos[15705]=-71;
cos[15706]=-71;
cos[15707]=-71;
cos[15708]=-71;
cos[15709]=-71;
cos[15710]=-70;
cos[15711]=-70;
cos[15712]=-70;
cos[15713]=-70;
cos[15714]=-70;
cos[15715]=-70;
cos[15716]=-70;
cos[15717]=-70;
cos[15718]=-70;
cos[15719]=-70;
cos[15720]=-70;
cos[15721]=-70;
cos[15722]=-70;
cos[15723]=-70;
cos[15724]=-70;
cos[15725]=-70;
cos[15726]=-70;
cos[15727]=-70;
cos[15728]=-70;
cos[15729]=-70;
cos[15730]=-70;
cos[15731]=-70;
cos[15732]=-70;
cos[15733]=-70;
cos[15734]=-70;
cos[15735]=-70;
cos[15736]=-70;
cos[15737]=-70;
cos[15738]=-70;
cos[15739]=-70;
cos[15740]=-70;
cos[15741]=-70;
cos[15742]=-70;
cos[15743]=-70;
cos[15744]=-70;
cos[15745]=-70;
cos[15746]=-70;
cos[15747]=-70;
cos[15748]=-70;
cos[15749]=-70;
cos[15750]=-70;
cos[15751]=-70;
cos[15752]=-70;
cos[15753]=-70;
cos[15754]=-70;
cos[15755]=-69;
cos[15756]=-69;
cos[15757]=-69;
cos[15758]=-69;
cos[15759]=-69;
cos[15760]=-69;
cos[15761]=-69;
cos[15762]=-69;
cos[15763]=-69;
cos[15764]=-69;
cos[15765]=-69;
cos[15766]=-69;
cos[15767]=-69;
cos[15768]=-69;
cos[15769]=-69;
cos[15770]=-69;
cos[15771]=-69;
cos[15772]=-69;
cos[15773]=-69;
cos[15774]=-69;
cos[15775]=-69;
cos[15776]=-69;
cos[15777]=-69;
cos[15778]=-69;
cos[15779]=-69;
cos[15780]=-69;
cos[15781]=-69;
cos[15782]=-69;
cos[15783]=-69;
cos[15784]=-69;
cos[15785]=-69;
cos[15786]=-69;
cos[15787]=-69;
cos[15788]=-69;
cos[15789]=-69;
cos[15790]=-69;
cos[15791]=-69;
cos[15792]=-69;
cos[15793]=-69;
cos[15794]=-69;
cos[15795]=-69;
cos[15796]=-69;
cos[15797]=-69;
cos[15798]=-69;
cos[15799]=-68;
cos[15800]=-68;
cos[15801]=-68;
cos[15802]=-68;
cos[15803]=-68;
cos[15804]=-68;
cos[15805]=-68;
cos[15806]=-68;
cos[15807]=-68;
cos[15808]=-68;
cos[15809]=-68;
cos[15810]=-68;
cos[15811]=-68;
cos[15812]=-68;
cos[15813]=-68;
cos[15814]=-68;
cos[15815]=-68;
cos[15816]=-68;
cos[15817]=-68;
cos[15818]=-68;
cos[15819]=-68;
cos[15820]=-68;
cos[15821]=-68;
cos[15822]=-68;
cos[15823]=-68;
cos[15824]=-68;
cos[15825]=-68;
cos[15826]=-68;
cos[15827]=-68;
cos[15828]=-68;
cos[15829]=-68;
cos[15830]=-68;
cos[15831]=-68;
cos[15832]=-68;
cos[15833]=-68;
cos[15834]=-68;
cos[15835]=-68;
cos[15836]=-68;
cos[15837]=-68;
cos[15838]=-68;
cos[15839]=-68;
cos[15840]=-67;
cos[15841]=-67;
cos[15842]=-67;
cos[15843]=-67;
cos[15844]=-67;
cos[15845]=-67;
cos[15846]=-67;
cos[15847]=-67;
cos[15848]=-67;
cos[15849]=-67;
cos[15850]=-67;
cos[15851]=-67;
cos[15852]=-67;
cos[15853]=-67;
cos[15854]=-67;
cos[15855]=-67;
cos[15856]=-67;
cos[15857]=-67;
cos[15858]=-67;
cos[15859]=-67;
cos[15860]=-67;
cos[15861]=-67;
cos[15862]=-67;
cos[15863]=-67;
cos[15864]=-67;
cos[15865]=-67;
cos[15866]=-67;
cos[15867]=-67;
cos[15868]=-67;
cos[15869]=-67;
cos[15870]=-67;
cos[15871]=-67;
cos[15872]=-67;
cos[15873]=-67;
cos[15874]=-67;
cos[15875]=-67;
cos[15876]=-67;
cos[15877]=-67;
cos[15878]=-67;
cos[15879]=-67;
cos[15880]=-66;
cos[15881]=-66;
cos[15882]=-66;
cos[15883]=-66;
cos[15884]=-66;
cos[15885]=-66;
cos[15886]=-66;
cos[15887]=-66;
cos[15888]=-66;
cos[15889]=-66;
cos[15890]=-66;
cos[15891]=-66;
cos[15892]=-66;
cos[15893]=-66;
cos[15894]=-66;
cos[15895]=-66;
cos[15896]=-66;
cos[15897]=-66;
cos[15898]=-66;
cos[15899]=-66;
cos[15900]=-66;
cos[15901]=-66;
cos[15902]=-66;
cos[15903]=-66;
cos[15904]=-66;
cos[15905]=-66;
cos[15906]=-66;
cos[15907]=-66;
cos[15908]=-66;
cos[15909]=-66;
cos[15910]=-66;
cos[15911]=-66;
cos[15912]=-66;
cos[15913]=-66;
cos[15914]=-66;
cos[15915]=-66;
cos[15916]=-66;
cos[15917]=-66;
cos[15918]=-65;
cos[15919]=-65;
cos[15920]=-65;
cos[15921]=-65;
cos[15922]=-65;
cos[15923]=-65;
cos[15924]=-65;
cos[15925]=-65;
cos[15926]=-65;
cos[15927]=-65;
cos[15928]=-65;
cos[15929]=-65;
cos[15930]=-65;
cos[15931]=-65;
cos[15932]=-65;
cos[15933]=-65;
cos[15934]=-65;
cos[15935]=-65;
cos[15936]=-65;
cos[15937]=-65;
cos[15938]=-65;
cos[15939]=-65;
cos[15940]=-65;
cos[15941]=-65;
cos[15942]=-65;
cos[15943]=-65;
cos[15944]=-65;
cos[15945]=-65;
cos[15946]=-65;
cos[15947]=-65;
cos[15948]=-65;
cos[15949]=-65;
cos[15950]=-65;
cos[15951]=-65;
cos[15952]=-65;
cos[15953]=-65;
cos[15954]=-65;
cos[15955]=-64;
cos[15956]=-64;
cos[15957]=-64;
cos[15958]=-64;
cos[15959]=-64;
cos[15960]=-64;
cos[15961]=-64;
cos[15962]=-64;
cos[15963]=-64;
cos[15964]=-64;
cos[15965]=-64;
cos[15966]=-64;
cos[15967]=-64;
cos[15968]=-64;
cos[15969]=-64;
cos[15970]=-64;
cos[15971]=-64;
cos[15972]=-64;
cos[15973]=-64;
cos[15974]=-64;
cos[15975]=-64;
cos[15976]=-64;
cos[15977]=-64;
cos[15978]=-64;
cos[15979]=-64;
cos[15980]=-64;
cos[15981]=-64;
cos[15982]=-64;
cos[15983]=-64;
cos[15984]=-64;
cos[15985]=-64;
cos[15986]=-64;
cos[15987]=-64;
cos[15988]=-64;
cos[15989]=-64;
cos[15990]=-63;
cos[15991]=-63;
cos[15992]=-63;
cos[15993]=-63;
cos[15994]=-63;
cos[15995]=-63;
cos[15996]=-63;
cos[15997]=-63;
cos[15998]=-63;
cos[15999]=-63;
cos[16000]=-63;
cos[16001]=-63;
cos[16002]=-63;
cos[16003]=-63;
cos[16004]=-63;
cos[16005]=-63;
cos[16006]=-63;
cos[16007]=-63;
cos[16008]=-63;
cos[16009]=-63;
cos[16010]=-63;
cos[16011]=-63;
cos[16012]=-63;
cos[16013]=-63;
cos[16014]=-63;
cos[16015]=-63;
cos[16016]=-63;
cos[16017]=-63;
cos[16018]=-63;
cos[16019]=-63;
cos[16020]=-63;
cos[16021]=-63;
cos[16022]=-63;
cos[16023]=-63;
cos[16024]=-63;
cos[16025]=-62;
cos[16026]=-62;
cos[16027]=-62;
cos[16028]=-62;
cos[16029]=-62;
cos[16030]=-62;
cos[16031]=-62;
cos[16032]=-62;
cos[16033]=-62;
cos[16034]=-62;
cos[16035]=-62;
cos[16036]=-62;
cos[16037]=-62;
cos[16038]=-62;
cos[16039]=-62;
cos[16040]=-62;
cos[16041]=-62;
cos[16042]=-62;
cos[16043]=-62;
cos[16044]=-62;
cos[16045]=-62;
cos[16046]=-62;
cos[16047]=-62;
cos[16048]=-62;
cos[16049]=-62;
cos[16050]=-62;
cos[16051]=-62;
cos[16052]=-62;
cos[16053]=-62;
cos[16054]=-62;
cos[16055]=-62;
cos[16056]=-62;
cos[16057]=-62;
cos[16058]=-61;
cos[16059]=-61;
cos[16060]=-61;
cos[16061]=-61;
cos[16062]=-61;
cos[16063]=-61;
cos[16064]=-61;
cos[16065]=-61;
cos[16066]=-61;
cos[16067]=-61;
cos[16068]=-61;
cos[16069]=-61;
cos[16070]=-61;
cos[16071]=-61;
cos[16072]=-61;
cos[16073]=-61;
cos[16074]=-61;
cos[16075]=-61;
cos[16076]=-61;
cos[16077]=-61;
cos[16078]=-61;
cos[16079]=-61;
cos[16080]=-61;
cos[16081]=-61;
cos[16082]=-61;
cos[16083]=-61;
cos[16084]=-61;
cos[16085]=-61;
cos[16086]=-61;
cos[16087]=-61;
cos[16088]=-61;
cos[16089]=-61;
cos[16090]=-61;
cos[16091]=-60;
cos[16092]=-60;
cos[16093]=-60;
cos[16094]=-60;
cos[16095]=-60;
cos[16096]=-60;
cos[16097]=-60;
cos[16098]=-60;
cos[16099]=-60;
cos[16100]=-60;
cos[16101]=-60;
cos[16102]=-60;
cos[16103]=-60;
cos[16104]=-60;
cos[16105]=-60;
cos[16106]=-60;
cos[16107]=-60;
cos[16108]=-60;
cos[16109]=-60;
cos[16110]=-60;
cos[16111]=-60;
cos[16112]=-60;
cos[16113]=-60;
cos[16114]=-60;
cos[16115]=-60;
cos[16116]=-60;
cos[16117]=-60;
cos[16118]=-60;
cos[16119]=-60;
cos[16120]=-60;
cos[16121]=-60;
cos[16122]=-60;
cos[16123]=-59;
cos[16124]=-59;
cos[16125]=-59;
cos[16126]=-59;
cos[16127]=-59;
cos[16128]=-59;
cos[16129]=-59;
cos[16130]=-59;
cos[16131]=-59;
cos[16132]=-59;
cos[16133]=-59;
cos[16134]=-59;
cos[16135]=-59;
cos[16136]=-59;
cos[16137]=-59;
cos[16138]=-59;
cos[16139]=-59;
cos[16140]=-59;
cos[16141]=-59;
cos[16142]=-59;
cos[16143]=-59;
cos[16144]=-59;
cos[16145]=-59;
cos[16146]=-59;
cos[16147]=-59;
cos[16148]=-59;
cos[16149]=-59;
cos[16150]=-59;
cos[16151]=-59;
cos[16152]=-59;
cos[16153]=-59;
cos[16154]=-58;
cos[16155]=-58;
cos[16156]=-58;
cos[16157]=-58;
cos[16158]=-58;
cos[16159]=-58;
cos[16160]=-58;
cos[16161]=-58;
cos[16162]=-58;
cos[16163]=-58;
cos[16164]=-58;
cos[16165]=-58;
cos[16166]=-58;
cos[16167]=-58;
cos[16168]=-58;
cos[16169]=-58;
cos[16170]=-58;
cos[16171]=-58;
cos[16172]=-58;
cos[16173]=-58;
cos[16174]=-58;
cos[16175]=-58;
cos[16176]=-58;
cos[16177]=-58;
cos[16178]=-58;
cos[16179]=-58;
cos[16180]=-58;
cos[16181]=-58;
cos[16182]=-58;
cos[16183]=-58;
cos[16184]=-57;
cos[16185]=-57;
cos[16186]=-57;
cos[16187]=-57;
cos[16188]=-57;
cos[16189]=-57;
cos[16190]=-57;
cos[16191]=-57;
cos[16192]=-57;
cos[16193]=-57;
cos[16194]=-57;
cos[16195]=-57;
cos[16196]=-57;
cos[16197]=-57;
cos[16198]=-57;
cos[16199]=-57;
cos[16200]=-57;
cos[16201]=-57;
cos[16202]=-57;
cos[16203]=-57;
cos[16204]=-57;
cos[16205]=-57;
cos[16206]=-57;
cos[16207]=-57;
cos[16208]=-57;
cos[16209]=-57;
cos[16210]=-57;
cos[16211]=-57;
cos[16212]=-57;
cos[16213]=-57;
cos[16214]=-56;
cos[16215]=-56;
cos[16216]=-56;
cos[16217]=-56;
cos[16218]=-56;
cos[16219]=-56;
cos[16220]=-56;
cos[16221]=-56;
cos[16222]=-56;
cos[16223]=-56;
cos[16224]=-56;
cos[16225]=-56;
cos[16226]=-56;
cos[16227]=-56;
cos[16228]=-56;
cos[16229]=-56;
cos[16230]=-56;
cos[16231]=-56;
cos[16232]=-56;
cos[16233]=-56;
cos[16234]=-56;
cos[16235]=-56;
cos[16236]=-56;
cos[16237]=-56;
cos[16238]=-56;
cos[16239]=-56;
cos[16240]=-56;
cos[16241]=-56;
cos[16242]=-56;
cos[16243]=-55;
cos[16244]=-55;
cos[16245]=-55;
cos[16246]=-55;
cos[16247]=-55;
cos[16248]=-55;
cos[16249]=-55;
cos[16250]=-55;
cos[16251]=-55;
cos[16252]=-55;
cos[16253]=-55;
cos[16254]=-55;
cos[16255]=-55;
cos[16256]=-55;
cos[16257]=-55;
cos[16258]=-55;
cos[16259]=-55;
cos[16260]=-55;
cos[16261]=-55;
cos[16262]=-55;
cos[16263]=-55;
cos[16264]=-55;
cos[16265]=-55;
cos[16266]=-55;
cos[16267]=-55;
cos[16268]=-55;
cos[16269]=-55;
cos[16270]=-55;
cos[16271]=-55;
cos[16272]=-54;
cos[16273]=-54;
cos[16274]=-54;
cos[16275]=-54;
cos[16276]=-54;
cos[16277]=-54;
cos[16278]=-54;
cos[16279]=-54;
cos[16280]=-54;
cos[16281]=-54;
cos[16282]=-54;
cos[16283]=-54;
cos[16284]=-54;
cos[16285]=-54;
cos[16286]=-54;
cos[16287]=-54;
cos[16288]=-54;
cos[16289]=-54;
cos[16290]=-54;
cos[16291]=-54;
cos[16292]=-54;
cos[16293]=-54;
cos[16294]=-54;
cos[16295]=-54;
cos[16296]=-54;
cos[16297]=-54;
cos[16298]=-54;
cos[16299]=-54;
cos[16300]=-53;
cos[16301]=-53;
cos[16302]=-53;
cos[16303]=-53;
cos[16304]=-53;
cos[16305]=-53;
cos[16306]=-53;
cos[16307]=-53;
cos[16308]=-53;
cos[16309]=-53;
cos[16310]=-53;
cos[16311]=-53;
cos[16312]=-53;
cos[16313]=-53;
cos[16314]=-53;
cos[16315]=-53;
cos[16316]=-53;
cos[16317]=-53;
cos[16318]=-53;
cos[16319]=-53;
cos[16320]=-53;
cos[16321]=-53;
cos[16322]=-53;
cos[16323]=-53;
cos[16324]=-53;
cos[16325]=-53;
cos[16326]=-53;
cos[16327]=-53;
cos[16328]=-52;
cos[16329]=-52;
cos[16330]=-52;
cos[16331]=-52;
cos[16332]=-52;
cos[16333]=-52;
cos[16334]=-52;
cos[16335]=-52;
cos[16336]=-52;
cos[16337]=-52;
cos[16338]=-52;
cos[16339]=-52;
cos[16340]=-52;
cos[16341]=-52;
cos[16342]=-52;
cos[16343]=-52;
cos[16344]=-52;
cos[16345]=-52;
cos[16346]=-52;
cos[16347]=-52;
cos[16348]=-52;
cos[16349]=-52;
cos[16350]=-52;
cos[16351]=-52;
cos[16352]=-52;
cos[16353]=-52;
cos[16354]=-52;
cos[16355]=-51;
cos[16356]=-51;
cos[16357]=-51;
cos[16358]=-51;
cos[16359]=-51;
cos[16360]=-51;
cos[16361]=-51;
cos[16362]=-51;
cos[16363]=-51;
cos[16364]=-51;
cos[16365]=-51;
cos[16366]=-51;
cos[16367]=-51;
cos[16368]=-51;
cos[16369]=-51;
cos[16370]=-51;
cos[16371]=-51;
cos[16372]=-51;
cos[16373]=-51;
cos[16374]=-51;
cos[16375]=-51;
cos[16376]=-51;
cos[16377]=-51;
cos[16378]=-51;
cos[16379]=-51;
cos[16380]=-51;
cos[16381]=-51;
cos[16382]=-50;
cos[16383]=-50;
cos[16384]=-50;
cos[16385]=-50;
cos[16386]=-50;
cos[16387]=-50;
cos[16388]=-50;
cos[16389]=-50;
cos[16390]=-50;
cos[16391]=-50;
cos[16392]=-50;
cos[16393]=-50;
cos[16394]=-50;
cos[16395]=-50;
cos[16396]=-50;
cos[16397]=-50;
cos[16398]=-50;
cos[16399]=-50;
cos[16400]=-50;
cos[16401]=-50;
cos[16402]=-50;
cos[16403]=-50;
cos[16404]=-50;
cos[16405]=-50;
cos[16406]=-50;
cos[16407]=-50;
cos[16408]=-49;
cos[16409]=-49;
cos[16410]=-49;
cos[16411]=-49;
cos[16412]=-49;
cos[16413]=-49;
cos[16414]=-49;
cos[16415]=-49;
cos[16416]=-49;
cos[16417]=-49;
cos[16418]=-49;
cos[16419]=-49;
cos[16420]=-49;
cos[16421]=-49;
cos[16422]=-49;
cos[16423]=-49;
cos[16424]=-49;
cos[16425]=-49;
cos[16426]=-49;
cos[16427]=-49;
cos[16428]=-49;
cos[16429]=-49;
cos[16430]=-49;
cos[16431]=-49;
cos[16432]=-49;
cos[16433]=-49;
cos[16434]=-49;
cos[16435]=-48;
cos[16436]=-48;
cos[16437]=-48;
cos[16438]=-48;
cos[16439]=-48;
cos[16440]=-48;
cos[16441]=-48;
cos[16442]=-48;
cos[16443]=-48;
cos[16444]=-48;
cos[16445]=-48;
cos[16446]=-48;
cos[16447]=-48;
cos[16448]=-48;
cos[16449]=-48;
cos[16450]=-48;
cos[16451]=-48;
cos[16452]=-48;
cos[16453]=-48;
cos[16454]=-48;
cos[16455]=-48;
cos[16456]=-48;
cos[16457]=-48;
cos[16458]=-48;
cos[16459]=-48;
cos[16460]=-47;
cos[16461]=-47;
cos[16462]=-47;
cos[16463]=-47;
cos[16464]=-47;
cos[16465]=-47;
cos[16466]=-47;
cos[16467]=-47;
cos[16468]=-47;
cos[16469]=-47;
cos[16470]=-47;
cos[16471]=-47;
cos[16472]=-47;
cos[16473]=-47;
cos[16474]=-47;
cos[16475]=-47;
cos[16476]=-47;
cos[16477]=-47;
cos[16478]=-47;
cos[16479]=-47;
cos[16480]=-47;
cos[16481]=-47;
cos[16482]=-47;
cos[16483]=-47;
cos[16484]=-47;
cos[16485]=-47;
cos[16486]=-46;
cos[16487]=-46;
cos[16488]=-46;
cos[16489]=-46;
cos[16490]=-46;
cos[16491]=-46;
cos[16492]=-46;
cos[16493]=-46;
cos[16494]=-46;
cos[16495]=-46;
cos[16496]=-46;
cos[16497]=-46;
cos[16498]=-46;
cos[16499]=-46;
cos[16500]=-46;
cos[16501]=-46;
cos[16502]=-46;
cos[16503]=-46;
cos[16504]=-46;
cos[16505]=-46;
cos[16506]=-46;
cos[16507]=-46;
cos[16508]=-46;
cos[16509]=-46;
cos[16510]=-46;
cos[16511]=-45;
cos[16512]=-45;
cos[16513]=-45;
cos[16514]=-45;
cos[16515]=-45;
cos[16516]=-45;
cos[16517]=-45;
cos[16518]=-45;
cos[16519]=-45;
cos[16520]=-45;
cos[16521]=-45;
cos[16522]=-45;
cos[16523]=-45;
cos[16524]=-45;
cos[16525]=-45;
cos[16526]=-45;
cos[16527]=-45;
cos[16528]=-45;
cos[16529]=-45;
cos[16530]=-45;
cos[16531]=-45;
cos[16532]=-45;
cos[16533]=-45;
cos[16534]=-45;
cos[16535]=-45;
cos[16536]=-44;
cos[16537]=-44;
cos[16538]=-44;
cos[16539]=-44;
cos[16540]=-44;
cos[16541]=-44;
cos[16542]=-44;
cos[16543]=-44;
cos[16544]=-44;
cos[16545]=-44;
cos[16546]=-44;
cos[16547]=-44;
cos[16548]=-44;
cos[16549]=-44;
cos[16550]=-44;
cos[16551]=-44;
cos[16552]=-44;
cos[16553]=-44;
cos[16554]=-44;
cos[16555]=-44;
cos[16556]=-44;
cos[16557]=-44;
cos[16558]=-44;
cos[16559]=-44;
cos[16560]=-44;
cos[16561]=-43;
cos[16562]=-43;
cos[16563]=-43;
cos[16564]=-43;
cos[16565]=-43;
cos[16566]=-43;
cos[16567]=-43;
cos[16568]=-43;
cos[16569]=-43;
cos[16570]=-43;
cos[16571]=-43;
cos[16572]=-43;
cos[16573]=-43;
cos[16574]=-43;
cos[16575]=-43;
cos[16576]=-43;
cos[16577]=-43;
cos[16578]=-43;
cos[16579]=-43;
cos[16580]=-43;
cos[16581]=-43;
cos[16582]=-43;
cos[16583]=-43;
cos[16584]=-43;
cos[16585]=-42;
cos[16586]=-42;
cos[16587]=-42;
cos[16588]=-42;
cos[16589]=-42;
cos[16590]=-42;
cos[16591]=-42;
cos[16592]=-42;
cos[16593]=-42;
cos[16594]=-42;
cos[16595]=-42;
cos[16596]=-42;
cos[16597]=-42;
cos[16598]=-42;
cos[16599]=-42;
cos[16600]=-42;
cos[16601]=-42;
cos[16602]=-42;
cos[16603]=-42;
cos[16604]=-42;
cos[16605]=-42;
cos[16606]=-42;
cos[16607]=-42;
cos[16608]=-42;
cos[16609]=-41;
cos[16610]=-41;
cos[16611]=-41;
cos[16612]=-41;
cos[16613]=-41;
cos[16614]=-41;
cos[16615]=-41;
cos[16616]=-41;
cos[16617]=-41;
cos[16618]=-41;
cos[16619]=-41;
cos[16620]=-41;
cos[16621]=-41;
cos[16622]=-41;
cos[16623]=-41;
cos[16624]=-41;
cos[16625]=-41;
cos[16626]=-41;
cos[16627]=-41;
cos[16628]=-41;
cos[16629]=-41;
cos[16630]=-41;
cos[16631]=-41;
cos[16632]=-41;
cos[16633]=-40;
cos[16634]=-40;
cos[16635]=-40;
cos[16636]=-40;
cos[16637]=-40;
cos[16638]=-40;
cos[16639]=-40;
cos[16640]=-40;
cos[16641]=-40;
cos[16642]=-40;
cos[16643]=-40;
cos[16644]=-40;
cos[16645]=-40;
cos[16646]=-40;
cos[16647]=-40;
cos[16648]=-40;
cos[16649]=-40;
cos[16650]=-40;
cos[16651]=-40;
cos[16652]=-40;
cos[16653]=-40;
cos[16654]=-40;
cos[16655]=-40;
cos[16656]=-40;
cos[16657]=-39;
cos[16658]=-39;
cos[16659]=-39;
cos[16660]=-39;
cos[16661]=-39;
cos[16662]=-39;
cos[16663]=-39;
cos[16664]=-39;
cos[16665]=-39;
cos[16666]=-39;
cos[16667]=-39;
cos[16668]=-39;
cos[16669]=-39;
cos[16670]=-39;
cos[16671]=-39;
cos[16672]=-39;
cos[16673]=-39;
cos[16674]=-39;
cos[16675]=-39;
cos[16676]=-39;
cos[16677]=-39;
cos[16678]=-39;
cos[16679]=-39;
cos[16680]=-38;
cos[16681]=-38;
cos[16682]=-38;
cos[16683]=-38;
cos[16684]=-38;
cos[16685]=-38;
cos[16686]=-38;
cos[16687]=-38;
cos[16688]=-38;
cos[16689]=-38;
cos[16690]=-38;
cos[16691]=-38;
cos[16692]=-38;
cos[16693]=-38;
cos[16694]=-38;
cos[16695]=-38;
cos[16696]=-38;
cos[16697]=-38;
cos[16698]=-38;
cos[16699]=-38;
cos[16700]=-38;
cos[16701]=-38;
cos[16702]=-38;
cos[16703]=-38;
cos[16704]=-37;
cos[16705]=-37;
cos[16706]=-37;
cos[16707]=-37;
cos[16708]=-37;
cos[16709]=-37;
cos[16710]=-37;
cos[16711]=-37;
cos[16712]=-37;
cos[16713]=-37;
cos[16714]=-37;
cos[16715]=-37;
cos[16716]=-37;
cos[16717]=-37;
cos[16718]=-37;
cos[16719]=-37;
cos[16720]=-37;
cos[16721]=-37;
cos[16722]=-37;
cos[16723]=-37;
cos[16724]=-37;
cos[16725]=-37;
cos[16726]=-37;
cos[16727]=-36;
cos[16728]=-36;
cos[16729]=-36;
cos[16730]=-36;
cos[16731]=-36;
cos[16732]=-36;
cos[16733]=-36;
cos[16734]=-36;
cos[16735]=-36;
cos[16736]=-36;
cos[16737]=-36;
cos[16738]=-36;
cos[16739]=-36;
cos[16740]=-36;
cos[16741]=-36;
cos[16742]=-36;
cos[16743]=-36;
cos[16744]=-36;
cos[16745]=-36;
cos[16746]=-36;
cos[16747]=-36;
cos[16748]=-36;
cos[16749]=-36;
cos[16750]=-35;
cos[16751]=-35;
cos[16752]=-35;
cos[16753]=-35;
cos[16754]=-35;
cos[16755]=-35;
cos[16756]=-35;
cos[16757]=-35;
cos[16758]=-35;
cos[16759]=-35;
cos[16760]=-35;
cos[16761]=-35;
cos[16762]=-35;
cos[16763]=-35;
cos[16764]=-35;
cos[16765]=-35;
cos[16766]=-35;
cos[16767]=-35;
cos[16768]=-35;
cos[16769]=-35;
cos[16770]=-35;
cos[16771]=-35;
cos[16772]=-35;
cos[16773]=-34;
cos[16774]=-34;
cos[16775]=-34;
cos[16776]=-34;
cos[16777]=-34;
cos[16778]=-34;
cos[16779]=-34;
cos[16780]=-34;
cos[16781]=-34;
cos[16782]=-34;
cos[16783]=-34;
cos[16784]=-34;
cos[16785]=-34;
cos[16786]=-34;
cos[16787]=-34;
cos[16788]=-34;
cos[16789]=-34;
cos[16790]=-34;
cos[16791]=-34;
cos[16792]=-34;
cos[16793]=-34;
cos[16794]=-34;
cos[16795]=-33;
cos[16796]=-33;
cos[16797]=-33;
cos[16798]=-33;
cos[16799]=-33;
cos[16800]=-33;
cos[16801]=-33;
cos[16802]=-33;
cos[16803]=-33;
cos[16804]=-33;
cos[16805]=-33;
cos[16806]=-33;
cos[16807]=-33;
cos[16808]=-33;
cos[16809]=-33;
cos[16810]=-33;
cos[16811]=-33;
cos[16812]=-33;
cos[16813]=-33;
cos[16814]=-33;
cos[16815]=-33;
cos[16816]=-33;
cos[16817]=-33;
cos[16818]=-32;
cos[16819]=-32;
cos[16820]=-32;
cos[16821]=-32;
cos[16822]=-32;
cos[16823]=-32;
cos[16824]=-32;
cos[16825]=-32;
cos[16826]=-32;
cos[16827]=-32;
cos[16828]=-32;
cos[16829]=-32;
cos[16830]=-32;
cos[16831]=-32;
cos[16832]=-32;
cos[16833]=-32;
cos[16834]=-32;
cos[16835]=-32;
cos[16836]=-32;
cos[16837]=-32;
cos[16838]=-32;
cos[16839]=-32;
cos[16840]=-31;
cos[16841]=-31;
cos[16842]=-31;
cos[16843]=-31;
cos[16844]=-31;
cos[16845]=-31;
cos[16846]=-31;
cos[16847]=-31;
cos[16848]=-31;
cos[16849]=-31;
cos[16850]=-31;
cos[16851]=-31;
cos[16852]=-31;
cos[16853]=-31;
cos[16854]=-31;
cos[16855]=-31;
cos[16856]=-31;
cos[16857]=-31;
cos[16858]=-31;
cos[16859]=-31;
cos[16860]=-31;
cos[16861]=-31;
cos[16862]=-30;
cos[16863]=-30;
cos[16864]=-30;
cos[16865]=-30;
cos[16866]=-30;
cos[16867]=-30;
cos[16868]=-30;
cos[16869]=-30;
cos[16870]=-30;
cos[16871]=-30;
cos[16872]=-30;
cos[16873]=-30;
cos[16874]=-30;
cos[16875]=-30;
cos[16876]=-30;
cos[16877]=-30;
cos[16878]=-30;
cos[16879]=-30;
cos[16880]=-30;
cos[16881]=-30;
cos[16882]=-30;
cos[16883]=-30;
cos[16884]=-29;
cos[16885]=-29;
cos[16886]=-29;
cos[16887]=-29;
cos[16888]=-29;
cos[16889]=-29;
cos[16890]=-29;
cos[16891]=-29;
cos[16892]=-29;
cos[16893]=-29;
cos[16894]=-29;
cos[16895]=-29;
cos[16896]=-29;
cos[16897]=-29;
cos[16898]=-29;
cos[16899]=-29;
cos[16900]=-29;
cos[16901]=-29;
cos[16902]=-29;
cos[16903]=-29;
cos[16904]=-29;
cos[16905]=-29;
cos[16906]=-28;
cos[16907]=-28;
cos[16908]=-28;
cos[16909]=-28;
cos[16910]=-28;
cos[16911]=-28;
cos[16912]=-28;
cos[16913]=-28;
cos[16914]=-28;
cos[16915]=-28;
cos[16916]=-28;
cos[16917]=-28;
cos[16918]=-28;
cos[16919]=-28;
cos[16920]=-28;
cos[16921]=-28;
cos[16922]=-28;
cos[16923]=-28;
cos[16924]=-28;
cos[16925]=-28;
cos[16926]=-28;
cos[16927]=-28;
cos[16928]=-27;
cos[16929]=-27;
cos[16930]=-27;
cos[16931]=-27;
cos[16932]=-27;
cos[16933]=-27;
cos[16934]=-27;
cos[16935]=-27;
cos[16936]=-27;
cos[16937]=-27;
cos[16938]=-27;
cos[16939]=-27;
cos[16940]=-27;
cos[16941]=-27;
cos[16942]=-27;
cos[16943]=-27;
cos[16944]=-27;
cos[16945]=-27;
cos[16946]=-27;
cos[16947]=-27;
cos[16948]=-27;
cos[16949]=-27;
cos[16950]=-26;
cos[16951]=-26;
cos[16952]=-26;
cos[16953]=-26;
cos[16954]=-26;
cos[16955]=-26;
cos[16956]=-26;
cos[16957]=-26;
cos[16958]=-26;
cos[16959]=-26;
cos[16960]=-26;
cos[16961]=-26;
cos[16962]=-26;
cos[16963]=-26;
cos[16964]=-26;
cos[16965]=-26;
cos[16966]=-26;
cos[16967]=-26;
cos[16968]=-26;
cos[16969]=-26;
cos[16970]=-26;
cos[16971]=-25;
cos[16972]=-25;
cos[16973]=-25;
cos[16974]=-25;
cos[16975]=-25;
cos[16976]=-25;
cos[16977]=-25;
cos[16978]=-25;
cos[16979]=-25;
cos[16980]=-25;
cos[16981]=-25;
cos[16982]=-25;
cos[16983]=-25;
cos[16984]=-25;
cos[16985]=-25;
cos[16986]=-25;
cos[16987]=-25;
cos[16988]=-25;
cos[16989]=-25;
cos[16990]=-25;
cos[16991]=-25;
cos[16992]=-25;
cos[16993]=-24;
cos[16994]=-24;
cos[16995]=-24;
cos[16996]=-24;
cos[16997]=-24;
cos[16998]=-24;
cos[16999]=-24;
cos[17000]=-24;
cos[17001]=-24;
cos[17002]=-24;
cos[17003]=-24;
cos[17004]=-24;
cos[17005]=-24;
cos[17006]=-24;
cos[17007]=-24;
cos[17008]=-24;
cos[17009]=-24;
cos[17010]=-24;
cos[17011]=-24;
cos[17012]=-24;
cos[17013]=-24;
cos[17014]=-23;
cos[17015]=-23;
cos[17016]=-23;
cos[17017]=-23;
cos[17018]=-23;
cos[17019]=-23;
cos[17020]=-23;
cos[17021]=-23;
cos[17022]=-23;
cos[17023]=-23;
cos[17024]=-23;
cos[17025]=-23;
cos[17026]=-23;
cos[17027]=-23;
cos[17028]=-23;
cos[17029]=-23;
cos[17030]=-23;
cos[17031]=-23;
cos[17032]=-23;
cos[17033]=-23;
cos[17034]=-23;
cos[17035]=-23;
cos[17036]=-22;
cos[17037]=-22;
cos[17038]=-22;
cos[17039]=-22;
cos[17040]=-22;
cos[17041]=-22;
cos[17042]=-22;
cos[17043]=-22;
cos[17044]=-22;
cos[17045]=-22;
cos[17046]=-22;
cos[17047]=-22;
cos[17048]=-22;
cos[17049]=-22;
cos[17050]=-22;
cos[17051]=-22;
cos[17052]=-22;
cos[17053]=-22;
cos[17054]=-22;
cos[17055]=-22;
cos[17056]=-22;
cos[17057]=-21;
cos[17058]=-21;
cos[17059]=-21;
cos[17060]=-21;
cos[17061]=-21;
cos[17062]=-21;
cos[17063]=-21;
cos[17064]=-21;
cos[17065]=-21;
cos[17066]=-21;
cos[17067]=-21;
cos[17068]=-21;
cos[17069]=-21;
cos[17070]=-21;
cos[17071]=-21;
cos[17072]=-21;
cos[17073]=-21;
cos[17074]=-21;
cos[17075]=-21;
cos[17076]=-21;
cos[17077]=-21;
cos[17078]=-20;
cos[17079]=-20;
cos[17080]=-20;
cos[17081]=-20;
cos[17082]=-20;
cos[17083]=-20;
cos[17084]=-20;
cos[17085]=-20;
cos[17086]=-20;
cos[17087]=-20;
cos[17088]=-20;
cos[17089]=-20;
cos[17090]=-20;
cos[17091]=-20;
cos[17092]=-20;
cos[17093]=-20;
cos[17094]=-20;
cos[17095]=-20;
cos[17096]=-20;
cos[17097]=-20;
cos[17098]=-20;
cos[17099]=-19;
cos[17100]=-19;
cos[17101]=-19;
cos[17102]=-19;
cos[17103]=-19;
cos[17104]=-19;
cos[17105]=-19;
cos[17106]=-19;
cos[17107]=-19;
cos[17108]=-19;
cos[17109]=-19;
cos[17110]=-19;
cos[17111]=-19;
cos[17112]=-19;
cos[17113]=-19;
cos[17114]=-19;
cos[17115]=-19;
cos[17116]=-19;
cos[17117]=-19;
cos[17118]=-19;
cos[17119]=-19;
cos[17120]=-18;
cos[17121]=-18;
cos[17122]=-18;
cos[17123]=-18;
cos[17124]=-18;
cos[17125]=-18;
cos[17126]=-18;
cos[17127]=-18;
cos[17128]=-18;
cos[17129]=-18;
cos[17130]=-18;
cos[17131]=-18;
cos[17132]=-18;
cos[17133]=-18;
cos[17134]=-18;
cos[17135]=-18;
cos[17136]=-18;
cos[17137]=-18;
cos[17138]=-18;
cos[17139]=-18;
cos[17140]=-18;
cos[17141]=-17;
cos[17142]=-17;
cos[17143]=-17;
cos[17144]=-17;
cos[17145]=-17;
cos[17146]=-17;
cos[17147]=-17;
cos[17148]=-17;
cos[17149]=-17;
cos[17150]=-17;
cos[17151]=-17;
cos[17152]=-17;
cos[17153]=-17;
cos[17154]=-17;
cos[17155]=-17;
cos[17156]=-17;
cos[17157]=-17;
cos[17158]=-17;
cos[17159]=-17;
cos[17160]=-17;
cos[17161]=-17;
cos[17162]=-16;
cos[17163]=-16;
cos[17164]=-16;
cos[17165]=-16;
cos[17166]=-16;
cos[17167]=-16;
cos[17168]=-16;
cos[17169]=-16;
cos[17170]=-16;
cos[17171]=-16;
cos[17172]=-16;
cos[17173]=-16;
cos[17174]=-16;
cos[17175]=-16;
cos[17176]=-16;
cos[17177]=-16;
cos[17178]=-16;
cos[17179]=-16;
cos[17180]=-16;
cos[17181]=-16;
cos[17182]=-16;
cos[17183]=-15;
cos[17184]=-15;
cos[17185]=-15;
cos[17186]=-15;
cos[17187]=-15;
cos[17188]=-15;
cos[17189]=-15;
cos[17190]=-15;
cos[17191]=-15;
cos[17192]=-15;
cos[17193]=-15;
cos[17194]=-15;
cos[17195]=-15;
cos[17196]=-15;
cos[17197]=-15;
cos[17198]=-15;
cos[17199]=-15;
cos[17200]=-15;
cos[17201]=-15;
cos[17202]=-15;
cos[17203]=-14;
cos[17204]=-14;
cos[17205]=-14;
cos[17206]=-14;
cos[17207]=-14;
cos[17208]=-14;
cos[17209]=-14;
cos[17210]=-14;
cos[17211]=-14;
cos[17212]=-14;
cos[17213]=-14;
cos[17214]=-14;
cos[17215]=-14;
cos[17216]=-14;
cos[17217]=-14;
cos[17218]=-14;
cos[17219]=-14;
cos[17220]=-14;
cos[17221]=-14;
cos[17222]=-14;
cos[17223]=-14;
cos[17224]=-13;
cos[17225]=-13;
cos[17226]=-13;
cos[17227]=-13;
cos[17228]=-13;
cos[17229]=-13;
cos[17230]=-13;
cos[17231]=-13;
cos[17232]=-13;
cos[17233]=-13;
cos[17234]=-13;
cos[17235]=-13;
cos[17236]=-13;
cos[17237]=-13;
cos[17238]=-13;
cos[17239]=-13;
cos[17240]=-13;
cos[17241]=-13;
cos[17242]=-13;
cos[17243]=-13;
cos[17244]=-13;
cos[17245]=-12;
cos[17246]=-12;
cos[17247]=-12;
cos[17248]=-12;
cos[17249]=-12;
cos[17250]=-12;
cos[17251]=-12;
cos[17252]=-12;
cos[17253]=-12;
cos[17254]=-12;
cos[17255]=-12;
cos[17256]=-12;
cos[17257]=-12;
cos[17258]=-12;
cos[17259]=-12;
cos[17260]=-12;
cos[17261]=-12;
cos[17262]=-12;
cos[17263]=-12;
cos[17264]=-12;
cos[17265]=-11;
cos[17266]=-11;
cos[17267]=-11;
cos[17268]=-11;
cos[17269]=-11;
cos[17270]=-11;
cos[17271]=-11;
cos[17272]=-11;
cos[17273]=-11;
cos[17274]=-11;
cos[17275]=-11;
cos[17276]=-11;
cos[17277]=-11;
cos[17278]=-11;
cos[17279]=-11;
cos[17280]=-11;
cos[17281]=-11;
cos[17282]=-11;
cos[17283]=-11;
cos[17284]=-11;
cos[17285]=-11;
cos[17286]=-10;
cos[17287]=-10;
cos[17288]=-10;
cos[17289]=-10;
cos[17290]=-10;
cos[17291]=-10;
cos[17292]=-10;
cos[17293]=-10;
cos[17294]=-10;
cos[17295]=-10;
cos[17296]=-10;
cos[17297]=-10;
cos[17298]=-10;
cos[17299]=-10;
cos[17300]=-10;
cos[17301]=-10;
cos[17302]=-10;
cos[17303]=-10;
cos[17304]=-10;
cos[17305]=-10;
cos[17306]=-9;
cos[17307]=-9;
cos[17308]=-9;
cos[17309]=-9;
cos[17310]=-9;
cos[17311]=-9;
cos[17312]=-9;
cos[17313]=-9;
cos[17314]=-9;
cos[17315]=-9;
cos[17316]=-9;
cos[17317]=-9;
cos[17318]=-9;
cos[17319]=-9;
cos[17320]=-9;
cos[17321]=-9;
cos[17322]=-9;
cos[17323]=-9;
cos[17324]=-9;
cos[17325]=-9;
cos[17326]=-9;
cos[17327]=-8;
cos[17328]=-8;
cos[17329]=-8;
cos[17330]=-8;
cos[17331]=-8;
cos[17332]=-8;
cos[17333]=-8;
cos[17334]=-8;
cos[17335]=-8;
cos[17336]=-8;
cos[17337]=-8;
cos[17338]=-8;
cos[17339]=-8;
cos[17340]=-8;
cos[17341]=-8;
cos[17342]=-8;
cos[17343]=-8;
cos[17344]=-8;
cos[17345]=-8;
cos[17346]=-8;
cos[17347]=-7;
cos[17348]=-7;
cos[17349]=-7;
cos[17350]=-7;
cos[17351]=-7;
cos[17352]=-7;
cos[17353]=-7;
cos[17354]=-7;
cos[17355]=-7;
cos[17356]=-7;
cos[17357]=-7;
cos[17358]=-7;
cos[17359]=-7;
cos[17360]=-7;
cos[17361]=-7;
cos[17362]=-7;
cos[17363]=-7;
cos[17364]=-7;
cos[17365]=-7;
cos[17366]=-7;
cos[17367]=-7;
cos[17368]=-6;
cos[17369]=-6;
cos[17370]=-6;
cos[17371]=-6;
cos[17372]=-6;
cos[17373]=-6;
cos[17374]=-6;
cos[17375]=-6;
cos[17376]=-6;
cos[17377]=-6;
cos[17378]=-6;
cos[17379]=-6;
cos[17380]=-6;
cos[17381]=-6;
cos[17382]=-6;
cos[17383]=-6;
cos[17384]=-6;
cos[17385]=-6;
cos[17386]=-6;
cos[17387]=-6;
cos[17388]=-5;
cos[17389]=-5;
cos[17390]=-5;
cos[17391]=-5;
cos[17392]=-5;
cos[17393]=-5;
cos[17394]=-5;
cos[17395]=-5;
cos[17396]=-5;
cos[17397]=-5;
cos[17398]=-5;
cos[17399]=-5;
cos[17400]=-5;
cos[17401]=-5;
cos[17402]=-5;
cos[17403]=-5;
cos[17404]=-5;
cos[17405]=-5;
cos[17406]=-5;
cos[17407]=-5;
cos[17408]=-5;
cos[17409]=-4;
cos[17410]=-4;
cos[17411]=-4;
cos[17412]=-4;
cos[17413]=-4;
cos[17414]=-4;
cos[17415]=-4;
cos[17416]=-4;
cos[17417]=-4;
cos[17418]=-4;
cos[17419]=-4;
cos[17420]=-4;
cos[17421]=-4;
cos[17422]=-4;
cos[17423]=-4;
cos[17424]=-4;
cos[17425]=-4;
cos[17426]=-4;
cos[17427]=-4;
cos[17428]=-4;
cos[17429]=-3;
cos[17430]=-3;
cos[17431]=-3;
cos[17432]=-3;
cos[17433]=-3;
cos[17434]=-3;
cos[17435]=-3;
cos[17436]=-3;
cos[17437]=-3;
cos[17438]=-3;
cos[17439]=-3;
cos[17440]=-3;
cos[17441]=-3;
cos[17442]=-3;
cos[17443]=-3;
cos[17444]=-3;
cos[17445]=-3;
cos[17446]=-3;
cos[17447]=-3;
cos[17448]=-3;
cos[17449]=-3;
cos[17450]=-2;
cos[17451]=-2;
cos[17452]=-2;
cos[17453]=-2;
cos[17454]=-2;
cos[17455]=-2;
cos[17456]=-2;
cos[17457]=-2;
cos[17458]=-2;
cos[17459]=-2;
cos[17460]=-2;
cos[17461]=-2;
cos[17462]=-2;
cos[17463]=-2;
cos[17464]=-2;
cos[17465]=-2;
cos[17466]=-2;
cos[17467]=-2;
cos[17468]=-2;
cos[17469]=-2;
cos[17470]=-1;
cos[17471]=-1;
cos[17472]=-1;
cos[17473]=-1;
cos[17474]=-1;
cos[17475]=-1;
cos[17476]=-1;
cos[17477]=-1;
cos[17478]=-1;
cos[17479]=-1;
cos[17480]=-1;
cos[17481]=-1;
cos[17482]=-1;
cos[17483]=-1;
cos[17484]=-1;
cos[17485]=-1;
cos[17486]=-1;
cos[17487]=-1;
cos[17488]=-1;
cos[17489]=-1;
cos[17490]=0;
cos[17491]=0;
cos[17492]=0;
cos[17493]=0;
cos[17494]=0;
cos[17495]=0;
cos[17496]=0;
cos[17497]=0;
cos[17498]=0;
cos[17499]=0;
cos[17500]=0;
cos[17501]=0;
cos[17502]=0;
cos[17503]=0;
cos[17504]=0;
cos[17505]=0;
cos[17506]=0;
cos[17507]=0;
cos[17508]=0;
cos[17509]=0;
cos[17510]=0;
cos[17511]=1;
cos[17512]=1;
cos[17513]=1;
cos[17514]=1;
cos[17515]=1;
cos[17516]=1;
cos[17517]=1;
cos[17518]=1;
cos[17519]=1;
cos[17520]=1;
cos[17521]=1;
cos[17522]=1;
cos[17523]=1;
cos[17524]=1;
cos[17525]=1;
cos[17526]=1;
cos[17527]=1;
cos[17528]=1;
cos[17529]=1;
cos[17530]=1;
cos[17531]=2;
cos[17532]=2;
cos[17533]=2;
cos[17534]=2;
cos[17535]=2;
cos[17536]=2;
cos[17537]=2;
cos[17538]=2;
cos[17539]=2;
cos[17540]=2;
cos[17541]=2;
cos[17542]=2;
cos[17543]=2;
cos[17544]=2;
cos[17545]=2;
cos[17546]=2;
cos[17547]=2;
cos[17548]=2;
cos[17549]=2;
cos[17550]=2;
cos[17551]=3;
cos[17552]=3;
cos[17553]=3;
cos[17554]=3;
cos[17555]=3;
cos[17556]=3;
cos[17557]=3;
cos[17558]=3;
cos[17559]=3;
cos[17560]=3;
cos[17561]=3;
cos[17562]=3;
cos[17563]=3;
cos[17564]=3;
cos[17565]=3;
cos[17566]=3;
cos[17567]=3;
cos[17568]=3;
cos[17569]=3;
cos[17570]=3;
cos[17571]=3;
cos[17572]=4;
cos[17573]=4;
cos[17574]=4;
cos[17575]=4;
cos[17576]=4;
cos[17577]=4;
cos[17578]=4;
cos[17579]=4;
cos[17580]=4;
cos[17581]=4;
cos[17582]=4;
cos[17583]=4;
cos[17584]=4;
cos[17585]=4;
cos[17586]=4;
cos[17587]=4;
cos[17588]=4;
cos[17589]=4;
cos[17590]=4;
cos[17591]=4;
cos[17592]=5;
cos[17593]=5;
cos[17594]=5;
cos[17595]=5;
cos[17596]=5;
cos[17597]=5;
cos[17598]=5;
cos[17599]=5;
cos[17600]=5;
cos[17601]=5;
cos[17602]=5;
cos[17603]=5;
cos[17604]=5;
cos[17605]=5;
cos[17606]=5;
cos[17607]=5;
cos[17608]=5;
cos[17609]=5;
cos[17610]=5;
cos[17611]=5;
cos[17612]=5;
cos[17613]=6;
cos[17614]=6;
cos[17615]=6;
cos[17616]=6;
cos[17617]=6;
cos[17618]=6;
cos[17619]=6;
cos[17620]=6;
cos[17621]=6;
cos[17622]=6;
cos[17623]=6;
cos[17624]=6;
cos[17625]=6;
cos[17626]=6;
cos[17627]=6;
cos[17628]=6;
cos[17629]=6;
cos[17630]=6;
cos[17631]=6;
cos[17632]=6;
cos[17633]=7;
cos[17634]=7;
cos[17635]=7;
cos[17636]=7;
cos[17637]=7;
cos[17638]=7;
cos[17639]=7;
cos[17640]=7;
cos[17641]=7;
cos[17642]=7;
cos[17643]=7;
cos[17644]=7;
cos[17645]=7;
cos[17646]=7;
cos[17647]=7;
cos[17648]=7;
cos[17649]=7;
cos[17650]=7;
cos[17651]=7;
cos[17652]=7;
cos[17653]=7;
cos[17654]=8;
cos[17655]=8;
cos[17656]=8;
cos[17657]=8;
cos[17658]=8;
cos[17659]=8;
cos[17660]=8;
cos[17661]=8;
cos[17662]=8;
cos[17663]=8;
cos[17664]=8;
cos[17665]=8;
cos[17666]=8;
cos[17667]=8;
cos[17668]=8;
cos[17669]=8;
cos[17670]=8;
cos[17671]=8;
cos[17672]=8;
cos[17673]=8;
cos[17674]=9;
cos[17675]=9;
cos[17676]=9;
cos[17677]=9;
cos[17678]=9;
cos[17679]=9;
cos[17680]=9;
cos[17681]=9;
cos[17682]=9;
cos[17683]=9;
cos[17684]=9;
cos[17685]=9;
cos[17686]=9;
cos[17687]=9;
cos[17688]=9;
cos[17689]=9;
cos[17690]=9;
cos[17691]=9;
cos[17692]=9;
cos[17693]=9;
cos[17694]=9;
cos[17695]=10;
cos[17696]=10;
cos[17697]=10;
cos[17698]=10;
cos[17699]=10;
cos[17700]=10;
cos[17701]=10;
cos[17702]=10;
cos[17703]=10;
cos[17704]=10;
cos[17705]=10;
cos[17706]=10;
cos[17707]=10;
cos[17708]=10;
cos[17709]=10;
cos[17710]=10;
cos[17711]=10;
cos[17712]=10;
cos[17713]=10;
cos[17714]=10;
cos[17715]=11;
cos[17716]=11;
cos[17717]=11;
cos[17718]=11;
cos[17719]=11;
cos[17720]=11;
cos[17721]=11;
cos[17722]=11;
cos[17723]=11;
cos[17724]=11;
cos[17725]=11;
cos[17726]=11;
cos[17727]=11;
cos[17728]=11;
cos[17729]=11;
cos[17730]=11;
cos[17731]=11;
cos[17732]=11;
cos[17733]=11;
cos[17734]=11;
cos[17735]=11;
cos[17736]=12;
cos[17737]=12;
cos[17738]=12;
cos[17739]=12;
cos[17740]=12;
cos[17741]=12;
cos[17742]=12;
cos[17743]=12;
cos[17744]=12;
cos[17745]=12;
cos[17746]=12;
cos[17747]=12;
cos[17748]=12;
cos[17749]=12;
cos[17750]=12;
cos[17751]=12;
cos[17752]=12;
cos[17753]=12;
cos[17754]=12;
cos[17755]=12;
cos[17756]=13;
cos[17757]=13;
cos[17758]=13;
cos[17759]=13;
cos[17760]=13;
cos[17761]=13;
cos[17762]=13;
cos[17763]=13;
cos[17764]=13;
cos[17765]=13;
cos[17766]=13;
cos[17767]=13;
cos[17768]=13;
cos[17769]=13;
cos[17770]=13;
cos[17771]=13;
cos[17772]=13;
cos[17773]=13;
cos[17774]=13;
cos[17775]=13;
cos[17776]=13;
cos[17777]=14;
cos[17778]=14;
cos[17779]=14;
cos[17780]=14;
cos[17781]=14;
cos[17782]=14;
cos[17783]=14;
cos[17784]=14;
cos[17785]=14;
cos[17786]=14;
cos[17787]=14;
cos[17788]=14;
cos[17789]=14;
cos[17790]=14;
cos[17791]=14;
cos[17792]=14;
cos[17793]=14;
cos[17794]=14;
cos[17795]=14;
cos[17796]=14;
cos[17797]=14;
cos[17798]=15;
cos[17799]=15;
cos[17800]=15;
cos[17801]=15;
cos[17802]=15;
cos[17803]=15;
cos[17804]=15;
cos[17805]=15;
cos[17806]=15;
cos[17807]=15;
cos[17808]=15;
cos[17809]=15;
cos[17810]=15;
cos[17811]=15;
cos[17812]=15;
cos[17813]=15;
cos[17814]=15;
cos[17815]=15;
cos[17816]=15;
cos[17817]=15;
cos[17818]=16;
cos[17819]=16;
cos[17820]=16;
cos[17821]=16;
cos[17822]=16;
cos[17823]=16;
cos[17824]=16;
cos[17825]=16;
cos[17826]=16;
cos[17827]=16;
cos[17828]=16;
cos[17829]=16;
cos[17830]=16;
cos[17831]=16;
cos[17832]=16;
cos[17833]=16;
cos[17834]=16;
cos[17835]=16;
cos[17836]=16;
cos[17837]=16;
cos[17838]=16;
cos[17839]=17;
cos[17840]=17;
cos[17841]=17;
cos[17842]=17;
cos[17843]=17;
cos[17844]=17;
cos[17845]=17;
cos[17846]=17;
cos[17847]=17;
cos[17848]=17;
cos[17849]=17;
cos[17850]=17;
cos[17851]=17;
cos[17852]=17;
cos[17853]=17;
cos[17854]=17;
cos[17855]=17;
cos[17856]=17;
cos[17857]=17;
cos[17858]=17;
cos[17859]=17;
cos[17860]=18;
cos[17861]=18;
cos[17862]=18;
cos[17863]=18;
cos[17864]=18;
cos[17865]=18;
cos[17866]=18;
cos[17867]=18;
cos[17868]=18;
cos[17869]=18;
cos[17870]=18;
cos[17871]=18;
cos[17872]=18;
cos[17873]=18;
cos[17874]=18;
cos[17875]=18;
cos[17876]=18;
cos[17877]=18;
cos[17878]=18;
cos[17879]=18;
cos[17880]=18;
cos[17881]=19;
cos[17882]=19;
cos[17883]=19;
cos[17884]=19;
cos[17885]=19;
cos[17886]=19;
cos[17887]=19;
cos[17888]=19;
cos[17889]=19;
cos[17890]=19;
cos[17891]=19;
cos[17892]=19;
cos[17893]=19;
cos[17894]=19;
cos[17895]=19;
cos[17896]=19;
cos[17897]=19;
cos[17898]=19;
cos[17899]=19;
cos[17900]=19;
cos[17901]=19;
cos[17902]=20;
cos[17903]=20;
cos[17904]=20;
cos[17905]=20;
cos[17906]=20;
cos[17907]=20;
cos[17908]=20;
cos[17909]=20;
cos[17910]=20;
cos[17911]=20;
cos[17912]=20;
cos[17913]=20;
cos[17914]=20;
cos[17915]=20;
cos[17916]=20;
cos[17917]=20;
cos[17918]=20;
cos[17919]=20;
cos[17920]=20;
cos[17921]=20;
cos[17922]=20;
cos[17923]=21;
cos[17924]=21;
cos[17925]=21;
cos[17926]=21;
cos[17927]=21;
cos[17928]=21;
cos[17929]=21;
cos[17930]=21;
cos[17931]=21;
cos[17932]=21;
cos[17933]=21;
cos[17934]=21;
cos[17935]=21;
cos[17936]=21;
cos[17937]=21;
cos[17938]=21;
cos[17939]=21;
cos[17940]=21;
cos[17941]=21;
cos[17942]=21;
cos[17943]=21;
cos[17944]=22;
cos[17945]=22;
cos[17946]=22;
cos[17947]=22;
cos[17948]=22;
cos[17949]=22;
cos[17950]=22;
cos[17951]=22;
cos[17952]=22;
cos[17953]=22;
cos[17954]=22;
cos[17955]=22;
cos[17956]=22;
cos[17957]=22;
cos[17958]=22;
cos[17959]=22;
cos[17960]=22;
cos[17961]=22;
cos[17962]=22;
cos[17963]=22;
cos[17964]=22;
cos[17965]=23;
cos[17966]=23;
cos[17967]=23;
cos[17968]=23;
cos[17969]=23;
cos[17970]=23;
cos[17971]=23;
cos[17972]=23;
cos[17973]=23;
cos[17974]=23;
cos[17975]=23;
cos[17976]=23;
cos[17977]=23;
cos[17978]=23;
cos[17979]=23;
cos[17980]=23;
cos[17981]=23;
cos[17982]=23;
cos[17983]=23;
cos[17984]=23;
cos[17985]=23;
cos[17986]=23;
cos[17987]=24;
cos[17988]=24;
cos[17989]=24;
cos[17990]=24;
cos[17991]=24;
cos[17992]=24;
cos[17993]=24;
cos[17994]=24;
cos[17995]=24;
cos[17996]=24;
cos[17997]=24;
cos[17998]=24;
cos[17999]=24;
cos[18000]=24;
cos[18001]=24;
cos[18002]=24;
cos[18003]=24;
cos[18004]=24;
cos[18005]=24;
cos[18006]=24;
cos[18007]=24;
cos[18008]=25;
cos[18009]=25;
cos[18010]=25;
cos[18011]=25;
cos[18012]=25;
cos[18013]=25;
cos[18014]=25;
cos[18015]=25;
cos[18016]=25;
cos[18017]=25;
cos[18018]=25;
cos[18019]=25;
cos[18020]=25;
cos[18021]=25;
cos[18022]=25;
cos[18023]=25;
cos[18024]=25;
cos[18025]=25;
cos[18026]=25;
cos[18027]=25;
cos[18028]=25;
cos[18029]=25;
cos[18030]=26;
cos[18031]=26;
cos[18032]=26;
cos[18033]=26;
cos[18034]=26;
cos[18035]=26;
cos[18036]=26;
cos[18037]=26;
cos[18038]=26;
cos[18039]=26;
cos[18040]=26;
cos[18041]=26;
cos[18042]=26;
cos[18043]=26;
cos[18044]=26;
cos[18045]=26;
cos[18046]=26;
cos[18047]=26;
cos[18048]=26;
cos[18049]=26;
cos[18050]=26;
cos[18051]=27;
cos[18052]=27;
cos[18053]=27;
cos[18054]=27;
cos[18055]=27;
cos[18056]=27;
cos[18057]=27;
cos[18058]=27;
cos[18059]=27;
cos[18060]=27;
cos[18061]=27;
cos[18062]=27;
cos[18063]=27;
cos[18064]=27;
cos[18065]=27;
cos[18066]=27;
cos[18067]=27;
cos[18068]=27;
cos[18069]=27;
cos[18070]=27;
cos[18071]=27;
cos[18072]=27;
cos[18073]=28;
cos[18074]=28;
cos[18075]=28;
cos[18076]=28;
cos[18077]=28;
cos[18078]=28;
cos[18079]=28;
cos[18080]=28;
cos[18081]=28;
cos[18082]=28;
cos[18083]=28;
cos[18084]=28;
cos[18085]=28;
cos[18086]=28;
cos[18087]=28;
cos[18088]=28;
cos[18089]=28;
cos[18090]=28;
cos[18091]=28;
cos[18092]=28;
cos[18093]=28;
cos[18094]=28;
cos[18095]=29;
cos[18096]=29;
cos[18097]=29;
cos[18098]=29;
cos[18099]=29;
cos[18100]=29;
cos[18101]=29;
cos[18102]=29;
cos[18103]=29;
cos[18104]=29;
cos[18105]=29;
cos[18106]=29;
cos[18107]=29;
cos[18108]=29;
cos[18109]=29;
cos[18110]=29;
cos[18111]=29;
cos[18112]=29;
cos[18113]=29;
cos[18114]=29;
cos[18115]=29;
cos[18116]=29;
cos[18117]=30;
cos[18118]=30;
cos[18119]=30;
cos[18120]=30;
cos[18121]=30;
cos[18122]=30;
cos[18123]=30;
cos[18124]=30;
cos[18125]=30;
cos[18126]=30;
cos[18127]=30;
cos[18128]=30;
cos[18129]=30;
cos[18130]=30;
cos[18131]=30;
cos[18132]=30;
cos[18133]=30;
cos[18134]=30;
cos[18135]=30;
cos[18136]=30;
cos[18137]=30;
cos[18138]=30;
cos[18139]=31;
cos[18140]=31;
cos[18141]=31;
cos[18142]=31;
cos[18143]=31;
cos[18144]=31;
cos[18145]=31;
cos[18146]=31;
cos[18147]=31;
cos[18148]=31;
cos[18149]=31;
cos[18150]=31;
cos[18151]=31;
cos[18152]=31;
cos[18153]=31;
cos[18154]=31;
cos[18155]=31;
cos[18156]=31;
cos[18157]=31;
cos[18158]=31;
cos[18159]=31;
cos[18160]=31;
cos[18161]=32;
cos[18162]=32;
cos[18163]=32;
cos[18164]=32;
cos[18165]=32;
cos[18166]=32;
cos[18167]=32;
cos[18168]=32;
cos[18169]=32;
cos[18170]=32;
cos[18171]=32;
cos[18172]=32;
cos[18173]=32;
cos[18174]=32;
cos[18175]=32;
cos[18176]=32;
cos[18177]=32;
cos[18178]=32;
cos[18179]=32;
cos[18180]=32;
cos[18181]=32;
cos[18182]=32;
cos[18183]=33;
cos[18184]=33;
cos[18185]=33;
cos[18186]=33;
cos[18187]=33;
cos[18188]=33;
cos[18189]=33;
cos[18190]=33;
cos[18191]=33;
cos[18192]=33;
cos[18193]=33;
cos[18194]=33;
cos[18195]=33;
cos[18196]=33;
cos[18197]=33;
cos[18198]=33;
cos[18199]=33;
cos[18200]=33;
cos[18201]=33;
cos[18202]=33;
cos[18203]=33;
cos[18204]=33;
cos[18205]=33;
cos[18206]=34;
cos[18207]=34;
cos[18208]=34;
cos[18209]=34;
cos[18210]=34;
cos[18211]=34;
cos[18212]=34;
cos[18213]=34;
cos[18214]=34;
cos[18215]=34;
cos[18216]=34;
cos[18217]=34;
cos[18218]=34;
cos[18219]=34;
cos[18220]=34;
cos[18221]=34;
cos[18222]=34;
cos[18223]=34;
cos[18224]=34;
cos[18225]=34;
cos[18226]=34;
cos[18227]=34;
cos[18228]=35;
cos[18229]=35;
cos[18230]=35;
cos[18231]=35;
cos[18232]=35;
cos[18233]=35;
cos[18234]=35;
cos[18235]=35;
cos[18236]=35;
cos[18237]=35;
cos[18238]=35;
cos[18239]=35;
cos[18240]=35;
cos[18241]=35;
cos[18242]=35;
cos[18243]=35;
cos[18244]=35;
cos[18245]=35;
cos[18246]=35;
cos[18247]=35;
cos[18248]=35;
cos[18249]=35;
cos[18250]=35;
cos[18251]=36;
cos[18252]=36;
cos[18253]=36;
cos[18254]=36;
cos[18255]=36;
cos[18256]=36;
cos[18257]=36;
cos[18258]=36;
cos[18259]=36;
cos[18260]=36;
cos[18261]=36;
cos[18262]=36;
cos[18263]=36;
cos[18264]=36;
cos[18265]=36;
cos[18266]=36;
cos[18267]=36;
cos[18268]=36;
cos[18269]=36;
cos[18270]=36;
cos[18271]=36;
cos[18272]=36;
cos[18273]=36;
cos[18274]=37;
cos[18275]=37;
cos[18276]=37;
cos[18277]=37;
cos[18278]=37;
cos[18279]=37;
cos[18280]=37;
cos[18281]=37;
cos[18282]=37;
cos[18283]=37;
cos[18284]=37;
cos[18285]=37;
cos[18286]=37;
cos[18287]=37;
cos[18288]=37;
cos[18289]=37;
cos[18290]=37;
cos[18291]=37;
cos[18292]=37;
cos[18293]=37;
cos[18294]=37;
cos[18295]=37;
cos[18296]=37;
cos[18297]=38;
cos[18298]=38;
cos[18299]=38;
cos[18300]=38;
cos[18301]=38;
cos[18302]=38;
cos[18303]=38;
cos[18304]=38;
cos[18305]=38;
cos[18306]=38;
cos[18307]=38;
cos[18308]=38;
cos[18309]=38;
cos[18310]=38;
cos[18311]=38;
cos[18312]=38;
cos[18313]=38;
cos[18314]=38;
cos[18315]=38;
cos[18316]=38;
cos[18317]=38;
cos[18318]=38;
cos[18319]=38;
cos[18320]=38;
cos[18321]=39;
cos[18322]=39;
cos[18323]=39;
cos[18324]=39;
cos[18325]=39;
cos[18326]=39;
cos[18327]=39;
cos[18328]=39;
cos[18329]=39;
cos[18330]=39;
cos[18331]=39;
cos[18332]=39;
cos[18333]=39;
cos[18334]=39;
cos[18335]=39;
cos[18336]=39;
cos[18337]=39;
cos[18338]=39;
cos[18339]=39;
cos[18340]=39;
cos[18341]=39;
cos[18342]=39;
cos[18343]=39;
cos[18344]=40;
cos[18345]=40;
cos[18346]=40;
cos[18347]=40;
cos[18348]=40;
cos[18349]=40;
cos[18350]=40;
cos[18351]=40;
cos[18352]=40;
cos[18353]=40;
cos[18354]=40;
cos[18355]=40;
cos[18356]=40;
cos[18357]=40;
cos[18358]=40;
cos[18359]=40;
cos[18360]=40;
cos[18361]=40;
cos[18362]=40;
cos[18363]=40;
cos[18364]=40;
cos[18365]=40;
cos[18366]=40;
cos[18367]=40;
cos[18368]=41;
cos[18369]=41;
cos[18370]=41;
cos[18371]=41;
cos[18372]=41;
cos[18373]=41;
cos[18374]=41;
cos[18375]=41;
cos[18376]=41;
cos[18377]=41;
cos[18378]=41;
cos[18379]=41;
cos[18380]=41;
cos[18381]=41;
cos[18382]=41;
cos[18383]=41;
cos[18384]=41;
cos[18385]=41;
cos[18386]=41;
cos[18387]=41;
cos[18388]=41;
cos[18389]=41;
cos[18390]=41;
cos[18391]=41;
cos[18392]=42;
cos[18393]=42;
cos[18394]=42;
cos[18395]=42;
cos[18396]=42;
cos[18397]=42;
cos[18398]=42;
cos[18399]=42;
cos[18400]=42;
cos[18401]=42;
cos[18402]=42;
cos[18403]=42;
cos[18404]=42;
cos[18405]=42;
cos[18406]=42;
cos[18407]=42;
cos[18408]=42;
cos[18409]=42;
cos[18410]=42;
cos[18411]=42;
cos[18412]=42;
cos[18413]=42;
cos[18414]=42;
cos[18415]=42;
cos[18416]=43;
cos[18417]=43;
cos[18418]=43;
cos[18419]=43;
cos[18420]=43;
cos[18421]=43;
cos[18422]=43;
cos[18423]=43;
cos[18424]=43;
cos[18425]=43;
cos[18426]=43;
cos[18427]=43;
cos[18428]=43;
cos[18429]=43;
cos[18430]=43;
cos[18431]=43;
cos[18432]=43;
cos[18433]=43;
cos[18434]=43;
cos[18435]=43;
cos[18436]=43;
cos[18437]=43;
cos[18438]=43;
cos[18439]=43;
cos[18440]=44;
cos[18441]=44;
cos[18442]=44;
cos[18443]=44;
cos[18444]=44;
cos[18445]=44;
cos[18446]=44;
cos[18447]=44;
cos[18448]=44;
cos[18449]=44;
cos[18450]=44;
cos[18451]=44;
cos[18452]=44;
cos[18453]=44;
cos[18454]=44;
cos[18455]=44;
cos[18456]=44;
cos[18457]=44;
cos[18458]=44;
cos[18459]=44;
cos[18460]=44;
cos[18461]=44;
cos[18462]=44;
cos[18463]=44;
cos[18464]=44;
cos[18465]=45;
cos[18466]=45;
cos[18467]=45;
cos[18468]=45;
cos[18469]=45;
cos[18470]=45;
cos[18471]=45;
cos[18472]=45;
cos[18473]=45;
cos[18474]=45;
cos[18475]=45;
cos[18476]=45;
cos[18477]=45;
cos[18478]=45;
cos[18479]=45;
cos[18480]=45;
cos[18481]=45;
cos[18482]=45;
cos[18483]=45;
cos[18484]=45;
cos[18485]=45;
cos[18486]=45;
cos[18487]=45;
cos[18488]=45;
cos[18489]=45;
cos[18490]=46;
cos[18491]=46;
cos[18492]=46;
cos[18493]=46;
cos[18494]=46;
cos[18495]=46;
cos[18496]=46;
cos[18497]=46;
cos[18498]=46;
cos[18499]=46;
cos[18500]=46;
cos[18501]=46;
cos[18502]=46;
cos[18503]=46;
cos[18504]=46;
cos[18505]=46;
cos[18506]=46;
cos[18507]=46;
cos[18508]=46;
cos[18509]=46;
cos[18510]=46;
cos[18511]=46;
cos[18512]=46;
cos[18513]=46;
cos[18514]=46;
cos[18515]=47;
cos[18516]=47;
cos[18517]=47;
cos[18518]=47;
cos[18519]=47;
cos[18520]=47;
cos[18521]=47;
cos[18522]=47;
cos[18523]=47;
cos[18524]=47;
cos[18525]=47;
cos[18526]=47;
cos[18527]=47;
cos[18528]=47;
cos[18529]=47;
cos[18530]=47;
cos[18531]=47;
cos[18532]=47;
cos[18533]=47;
cos[18534]=47;
cos[18535]=47;
cos[18536]=47;
cos[18537]=47;
cos[18538]=47;
cos[18539]=47;
cos[18540]=47;
cos[18541]=48;
cos[18542]=48;
cos[18543]=48;
cos[18544]=48;
cos[18545]=48;
cos[18546]=48;
cos[18547]=48;
cos[18548]=48;
cos[18549]=48;
cos[18550]=48;
cos[18551]=48;
cos[18552]=48;
cos[18553]=48;
cos[18554]=48;
cos[18555]=48;
cos[18556]=48;
cos[18557]=48;
cos[18558]=48;
cos[18559]=48;
cos[18560]=48;
cos[18561]=48;
cos[18562]=48;
cos[18563]=48;
cos[18564]=48;
cos[18565]=48;
cos[18566]=49;
cos[18567]=49;
cos[18568]=49;
cos[18569]=49;
cos[18570]=49;
cos[18571]=49;
cos[18572]=49;
cos[18573]=49;
cos[18574]=49;
cos[18575]=49;
cos[18576]=49;
cos[18577]=49;
cos[18578]=49;
cos[18579]=49;
cos[18580]=49;
cos[18581]=49;
cos[18582]=49;
cos[18583]=49;
cos[18584]=49;
cos[18585]=49;
cos[18586]=49;
cos[18587]=49;
cos[18588]=49;
cos[18589]=49;
cos[18590]=49;
cos[18591]=49;
cos[18592]=49;
cos[18593]=50;
cos[18594]=50;
cos[18595]=50;
cos[18596]=50;
cos[18597]=50;
cos[18598]=50;
cos[18599]=50;
cos[18600]=50;
cos[18601]=50;
cos[18602]=50;
cos[18603]=50;
cos[18604]=50;
cos[18605]=50;
cos[18606]=50;
cos[18607]=50;
cos[18608]=50;
cos[18609]=50;
cos[18610]=50;
cos[18611]=50;
cos[18612]=50;
cos[18613]=50;
cos[18614]=50;
cos[18615]=50;
cos[18616]=50;
cos[18617]=50;
cos[18618]=50;
cos[18619]=51;
cos[18620]=51;
cos[18621]=51;
cos[18622]=51;
cos[18623]=51;
cos[18624]=51;
cos[18625]=51;
cos[18626]=51;
cos[18627]=51;
cos[18628]=51;
cos[18629]=51;
cos[18630]=51;
cos[18631]=51;
cos[18632]=51;
cos[18633]=51;
cos[18634]=51;
cos[18635]=51;
cos[18636]=51;
cos[18637]=51;
cos[18638]=51;
cos[18639]=51;
cos[18640]=51;
cos[18641]=51;
cos[18642]=51;
cos[18643]=51;
cos[18644]=51;
cos[18645]=51;
cos[18646]=52;
cos[18647]=52;
cos[18648]=52;
cos[18649]=52;
cos[18650]=52;
cos[18651]=52;
cos[18652]=52;
cos[18653]=52;
cos[18654]=52;
cos[18655]=52;
cos[18656]=52;
cos[18657]=52;
cos[18658]=52;
cos[18659]=52;
cos[18660]=52;
cos[18661]=52;
cos[18662]=52;
cos[18663]=52;
cos[18664]=52;
cos[18665]=52;
cos[18666]=52;
cos[18667]=52;
cos[18668]=52;
cos[18669]=52;
cos[18670]=52;
cos[18671]=52;
cos[18672]=52;
cos[18673]=53;
cos[18674]=53;
cos[18675]=53;
cos[18676]=53;
cos[18677]=53;
cos[18678]=53;
cos[18679]=53;
cos[18680]=53;
cos[18681]=53;
cos[18682]=53;
cos[18683]=53;
cos[18684]=53;
cos[18685]=53;
cos[18686]=53;
cos[18687]=53;
cos[18688]=53;
cos[18689]=53;
cos[18690]=53;
cos[18691]=53;
cos[18692]=53;
cos[18693]=53;
cos[18694]=53;
cos[18695]=53;
cos[18696]=53;
cos[18697]=53;
cos[18698]=53;
cos[18699]=53;
cos[18700]=53;
cos[18701]=54;
cos[18702]=54;
cos[18703]=54;
cos[18704]=54;
cos[18705]=54;
cos[18706]=54;
cos[18707]=54;
cos[18708]=54;
cos[18709]=54;
cos[18710]=54;
cos[18711]=54;
cos[18712]=54;
cos[18713]=54;
cos[18714]=54;
cos[18715]=54;
cos[18716]=54;
cos[18717]=54;
cos[18718]=54;
cos[18719]=54;
cos[18720]=54;
cos[18721]=54;
cos[18722]=54;
cos[18723]=54;
cos[18724]=54;
cos[18725]=54;
cos[18726]=54;
cos[18727]=54;
cos[18728]=54;
cos[18729]=55;
cos[18730]=55;
cos[18731]=55;
cos[18732]=55;
cos[18733]=55;
cos[18734]=55;
cos[18735]=55;
cos[18736]=55;
cos[18737]=55;
cos[18738]=55;
cos[18739]=55;
cos[18740]=55;
cos[18741]=55;
cos[18742]=55;
cos[18743]=55;
cos[18744]=55;
cos[18745]=55;
cos[18746]=55;
cos[18747]=55;
cos[18748]=55;
cos[18749]=55;
cos[18750]=55;
cos[18751]=55;
cos[18752]=55;
cos[18753]=55;
cos[18754]=55;
cos[18755]=55;
cos[18756]=55;
cos[18757]=55;
cos[18758]=56;
cos[18759]=56;
cos[18760]=56;
cos[18761]=56;
cos[18762]=56;
cos[18763]=56;
cos[18764]=56;
cos[18765]=56;
cos[18766]=56;
cos[18767]=56;
cos[18768]=56;
cos[18769]=56;
cos[18770]=56;
cos[18771]=56;
cos[18772]=56;
cos[18773]=56;
cos[18774]=56;
cos[18775]=56;
cos[18776]=56;
cos[18777]=56;
cos[18778]=56;
cos[18779]=56;
cos[18780]=56;
cos[18781]=56;
cos[18782]=56;
cos[18783]=56;
cos[18784]=56;
cos[18785]=56;
cos[18786]=56;
cos[18787]=57;
cos[18788]=57;
cos[18789]=57;
cos[18790]=57;
cos[18791]=57;
cos[18792]=57;
cos[18793]=57;
cos[18794]=57;
cos[18795]=57;
cos[18796]=57;
cos[18797]=57;
cos[18798]=57;
cos[18799]=57;
cos[18800]=57;
cos[18801]=57;
cos[18802]=57;
cos[18803]=57;
cos[18804]=57;
cos[18805]=57;
cos[18806]=57;
cos[18807]=57;
cos[18808]=57;
cos[18809]=57;
cos[18810]=57;
cos[18811]=57;
cos[18812]=57;
cos[18813]=57;
cos[18814]=57;
cos[18815]=57;
cos[18816]=57;
cos[18817]=58;
cos[18818]=58;
cos[18819]=58;
cos[18820]=58;
cos[18821]=58;
cos[18822]=58;
cos[18823]=58;
cos[18824]=58;
cos[18825]=58;
cos[18826]=58;
cos[18827]=58;
cos[18828]=58;
cos[18829]=58;
cos[18830]=58;
cos[18831]=58;
cos[18832]=58;
cos[18833]=58;
cos[18834]=58;
cos[18835]=58;
cos[18836]=58;
cos[18837]=58;
cos[18838]=58;
cos[18839]=58;
cos[18840]=58;
cos[18841]=58;
cos[18842]=58;
cos[18843]=58;
cos[18844]=58;
cos[18845]=58;
cos[18846]=58;
cos[18847]=59;
cos[18848]=59;
cos[18849]=59;
cos[18850]=59;
cos[18851]=59;
cos[18852]=59;
cos[18853]=59;
cos[18854]=59;
cos[18855]=59;
cos[18856]=59;
cos[18857]=59;
cos[18858]=59;
cos[18859]=59;
cos[18860]=59;
cos[18861]=59;
cos[18862]=59;
cos[18863]=59;
cos[18864]=59;
cos[18865]=59;
cos[18866]=59;
cos[18867]=59;
cos[18868]=59;
cos[18869]=59;
cos[18870]=59;
cos[18871]=59;
cos[18872]=59;
cos[18873]=59;
cos[18874]=59;
cos[18875]=59;
cos[18876]=59;
cos[18877]=59;
cos[18878]=60;
cos[18879]=60;
cos[18880]=60;
cos[18881]=60;
cos[18882]=60;
cos[18883]=60;
cos[18884]=60;
cos[18885]=60;
cos[18886]=60;
cos[18887]=60;
cos[18888]=60;
cos[18889]=60;
cos[18890]=60;
cos[18891]=60;
cos[18892]=60;
cos[18893]=60;
cos[18894]=60;
cos[18895]=60;
cos[18896]=60;
cos[18897]=60;
cos[18898]=60;
cos[18899]=60;
cos[18900]=60;
cos[18901]=60;
cos[18902]=60;
cos[18903]=60;
cos[18904]=60;
cos[18905]=60;
cos[18906]=60;
cos[18907]=60;
cos[18908]=60;
cos[18909]=60;
cos[18910]=61;
cos[18911]=61;
cos[18912]=61;
cos[18913]=61;
cos[18914]=61;
cos[18915]=61;
cos[18916]=61;
cos[18917]=61;
cos[18918]=61;
cos[18919]=61;
cos[18920]=61;
cos[18921]=61;
cos[18922]=61;
cos[18923]=61;
cos[18924]=61;
cos[18925]=61;
cos[18926]=61;
cos[18927]=61;
cos[18928]=61;
cos[18929]=61;
cos[18930]=61;
cos[18931]=61;
cos[18932]=61;
cos[18933]=61;
cos[18934]=61;
cos[18935]=61;
cos[18936]=61;
cos[18937]=61;
cos[18938]=61;
cos[18939]=61;
cos[18940]=61;
cos[18941]=61;
cos[18942]=61;
cos[18943]=62;
cos[18944]=62;
cos[18945]=62;
cos[18946]=62;
cos[18947]=62;
cos[18948]=62;
cos[18949]=62;
cos[18950]=62;
cos[18951]=62;
cos[18952]=62;
cos[18953]=62;
cos[18954]=62;
cos[18955]=62;
cos[18956]=62;
cos[18957]=62;
cos[18958]=62;
cos[18959]=62;
cos[18960]=62;
cos[18961]=62;
cos[18962]=62;
cos[18963]=62;
cos[18964]=62;
cos[18965]=62;
cos[18966]=62;
cos[18967]=62;
cos[18968]=62;
cos[18969]=62;
cos[18970]=62;
cos[18971]=62;
cos[18972]=62;
cos[18973]=62;
cos[18974]=62;
cos[18975]=62;
cos[18976]=63;
cos[18977]=63;
cos[18978]=63;
cos[18979]=63;
cos[18980]=63;
cos[18981]=63;
cos[18982]=63;
cos[18983]=63;
cos[18984]=63;
cos[18985]=63;
cos[18986]=63;
cos[18987]=63;
cos[18988]=63;
cos[18989]=63;
cos[18990]=63;
cos[18991]=63;
cos[18992]=63;
cos[18993]=63;
cos[18994]=63;
cos[18995]=63;
cos[18996]=63;
cos[18997]=63;
cos[18998]=63;
cos[18999]=63;
cos[19000]=63;
cos[19001]=63;
cos[19002]=63;
cos[19003]=63;
cos[19004]=63;
cos[19005]=63;
cos[19006]=63;
cos[19007]=63;
cos[19008]=63;
cos[19009]=63;
cos[19010]=63;
cos[19011]=64;
cos[19012]=64;
cos[19013]=64;
cos[19014]=64;
cos[19015]=64;
cos[19016]=64;
cos[19017]=64;
cos[19018]=64;
cos[19019]=64;
cos[19020]=64;
cos[19021]=64;
cos[19022]=64;
cos[19023]=64;
cos[19024]=64;
cos[19025]=64;
cos[19026]=64;
cos[19027]=64;
cos[19028]=64;
cos[19029]=64;
cos[19030]=64;
cos[19031]=64;
cos[19032]=64;
cos[19033]=64;
cos[19034]=64;
cos[19035]=64;
cos[19036]=64;
cos[19037]=64;
cos[19038]=64;
cos[19039]=64;
cos[19040]=64;
cos[19041]=64;
cos[19042]=64;
cos[19043]=64;
cos[19044]=64;
cos[19045]=64;
cos[19046]=65;
cos[19047]=65;
cos[19048]=65;
cos[19049]=65;
cos[19050]=65;
cos[19051]=65;
cos[19052]=65;
cos[19053]=65;
cos[19054]=65;
cos[19055]=65;
cos[19056]=65;
cos[19057]=65;
cos[19058]=65;
cos[19059]=65;
cos[19060]=65;
cos[19061]=65;
cos[19062]=65;
cos[19063]=65;
cos[19064]=65;
cos[19065]=65;
cos[19066]=65;
cos[19067]=65;
cos[19068]=65;
cos[19069]=65;
cos[19070]=65;
cos[19071]=65;
cos[19072]=65;
cos[19073]=65;
cos[19074]=65;
cos[19075]=65;
cos[19076]=65;
cos[19077]=65;
cos[19078]=65;
cos[19079]=65;
cos[19080]=65;
cos[19081]=65;
cos[19082]=65;
cos[19083]=66;
cos[19084]=66;
cos[19085]=66;
cos[19086]=66;
cos[19087]=66;
cos[19088]=66;
cos[19089]=66;
cos[19090]=66;
cos[19091]=66;
cos[19092]=66;
cos[19093]=66;
cos[19094]=66;
cos[19095]=66;
cos[19096]=66;
cos[19097]=66;
cos[19098]=66;
cos[19099]=66;
cos[19100]=66;
cos[19101]=66;
cos[19102]=66;
cos[19103]=66;
cos[19104]=66;
cos[19105]=66;
cos[19106]=66;
cos[19107]=66;
cos[19108]=66;
cos[19109]=66;
cos[19110]=66;
cos[19111]=66;
cos[19112]=66;
cos[19113]=66;
cos[19114]=66;
cos[19115]=66;
cos[19116]=66;
cos[19117]=66;
cos[19118]=66;
cos[19119]=66;
cos[19120]=66;
cos[19121]=67;
cos[19122]=67;
cos[19123]=67;
cos[19124]=67;
cos[19125]=67;
cos[19126]=67;
cos[19127]=67;
cos[19128]=67;
cos[19129]=67;
cos[19130]=67;
cos[19131]=67;
cos[19132]=67;
cos[19133]=67;
cos[19134]=67;
cos[19135]=67;
cos[19136]=67;
cos[19137]=67;
cos[19138]=67;
cos[19139]=67;
cos[19140]=67;
cos[19141]=67;
cos[19142]=67;
cos[19143]=67;
cos[19144]=67;
cos[19145]=67;
cos[19146]=67;
cos[19147]=67;
cos[19148]=67;
cos[19149]=67;
cos[19150]=67;
cos[19151]=67;
cos[19152]=67;
cos[19153]=67;
cos[19154]=67;
cos[19155]=67;
cos[19156]=67;
cos[19157]=67;
cos[19158]=67;
cos[19159]=67;
cos[19160]=67;
cos[19161]=68;
cos[19162]=68;
cos[19163]=68;
cos[19164]=68;
cos[19165]=68;
cos[19166]=68;
cos[19167]=68;
cos[19168]=68;
cos[19169]=68;
cos[19170]=68;
cos[19171]=68;
cos[19172]=68;
cos[19173]=68;
cos[19174]=68;
cos[19175]=68;
cos[19176]=68;
cos[19177]=68;
cos[19178]=68;
cos[19179]=68;
cos[19180]=68;
cos[19181]=68;
cos[19182]=68;
cos[19183]=68;
cos[19184]=68;
cos[19185]=68;
cos[19186]=68;
cos[19187]=68;
cos[19188]=68;
cos[19189]=68;
cos[19190]=68;
cos[19191]=68;
cos[19192]=68;
cos[19193]=68;
cos[19194]=68;
cos[19195]=68;
cos[19196]=68;
cos[19197]=68;
cos[19198]=68;
cos[19199]=68;
cos[19200]=68;
cos[19201]=68;
cos[19202]=69;
cos[19203]=69;
cos[19204]=69;
cos[19205]=69;
cos[19206]=69;
cos[19207]=69;
cos[19208]=69;
cos[19209]=69;
cos[19210]=69;
cos[19211]=69;
cos[19212]=69;
cos[19213]=69;
cos[19214]=69;
cos[19215]=69;
cos[19216]=69;
cos[19217]=69;
cos[19218]=69;
cos[19219]=69;
cos[19220]=69;
cos[19221]=69;
cos[19222]=69;
cos[19223]=69;
cos[19224]=69;
cos[19225]=69;
cos[19226]=69;
cos[19227]=69;
cos[19228]=69;
cos[19229]=69;
cos[19230]=69;
cos[19231]=69;
cos[19232]=69;
cos[19233]=69;
cos[19234]=69;
cos[19235]=69;
cos[19236]=69;
cos[19237]=69;
cos[19238]=69;
cos[19239]=69;
cos[19240]=69;
cos[19241]=69;
cos[19242]=69;
cos[19243]=69;
cos[19244]=69;
cos[19245]=69;
cos[19246]=70;
cos[19247]=70;
cos[19248]=70;
cos[19249]=70;
cos[19250]=70;
cos[19251]=70;
cos[19252]=70;
cos[19253]=70;
cos[19254]=70;
cos[19255]=70;
cos[19256]=70;
cos[19257]=70;
cos[19258]=70;
cos[19259]=70;
cos[19260]=70;
cos[19261]=70;
cos[19262]=70;
cos[19263]=70;
cos[19264]=70;
cos[19265]=70;
cos[19266]=70;
cos[19267]=70;
cos[19268]=70;
cos[19269]=70;
cos[19270]=70;
cos[19271]=70;
cos[19272]=70;
cos[19273]=70;
cos[19274]=70;
cos[19275]=70;
cos[19276]=70;
cos[19277]=70;
cos[19278]=70;
cos[19279]=70;
cos[19280]=70;
cos[19281]=70;
cos[19282]=70;
cos[19283]=70;
cos[19284]=70;
cos[19285]=70;
cos[19286]=70;
cos[19287]=70;
cos[19288]=70;
cos[19289]=70;
cos[19290]=70;
cos[19291]=71;
cos[19292]=71;
cos[19293]=71;
cos[19294]=71;
cos[19295]=71;
cos[19296]=71;
cos[19297]=71;
cos[19298]=71;
cos[19299]=71;
cos[19300]=71;
cos[19301]=71;
cos[19302]=71;
cos[19303]=71;
cos[19304]=71;
cos[19305]=71;
cos[19306]=71;
cos[19307]=71;
cos[19308]=71;
cos[19309]=71;
cos[19310]=71;
cos[19311]=71;
cos[19312]=71;
cos[19313]=71;
cos[19314]=71;
cos[19315]=71;
cos[19316]=71;
cos[19317]=71;
cos[19318]=71;
cos[19319]=71;
cos[19320]=71;
cos[19321]=71;
cos[19322]=71;
cos[19323]=71;
cos[19324]=71;
cos[19325]=71;
cos[19326]=71;
cos[19327]=71;
cos[19328]=71;
cos[19329]=71;
cos[19330]=71;
cos[19331]=71;
cos[19332]=71;
cos[19333]=71;
cos[19334]=71;
cos[19335]=71;
cos[19336]=71;
cos[19337]=71;
cos[19338]=71;
cos[19339]=71;
cos[19340]=72;
cos[19341]=72;
cos[19342]=72;
cos[19343]=72;
cos[19344]=72;
cos[19345]=72;
cos[19346]=72;
cos[19347]=72;
cos[19348]=72;
cos[19349]=72;
cos[19350]=72;
cos[19351]=72;
cos[19352]=72;
cos[19353]=72;
cos[19354]=72;
cos[19355]=72;
cos[19356]=72;
cos[19357]=72;
cos[19358]=72;
cos[19359]=72;
cos[19360]=72;
cos[19361]=72;
cos[19362]=72;
cos[19363]=72;
cos[19364]=72;
cos[19365]=72;
cos[19366]=72;
cos[19367]=72;
cos[19368]=72;
cos[19369]=72;
cos[19370]=72;
cos[19371]=72;
cos[19372]=72;
cos[19373]=72;
cos[19374]=72;
cos[19375]=72;
cos[19376]=72;
cos[19377]=72;
cos[19378]=72;
cos[19379]=72;
cos[19380]=72;
cos[19381]=72;
cos[19382]=72;
cos[19383]=72;
cos[19384]=72;
cos[19385]=72;
cos[19386]=72;
cos[19387]=72;
cos[19388]=72;
cos[19389]=72;
cos[19390]=72;
cos[19391]=72;
cos[19392]=72;
cos[19393]=73;
cos[19394]=73;
cos[19395]=73;
cos[19396]=73;
cos[19397]=73;
cos[19398]=73;
cos[19399]=73;
cos[19400]=73;
cos[19401]=73;
cos[19402]=73;
cos[19403]=73;
cos[19404]=73;
cos[19405]=73;
cos[19406]=73;
cos[19407]=73;
cos[19408]=73;
cos[19409]=73;
cos[19410]=73;
cos[19411]=73;
cos[19412]=73;
cos[19413]=73;
cos[19414]=73;
cos[19415]=73;
cos[19416]=73;
cos[19417]=73;
cos[19418]=73;
cos[19419]=73;
cos[19420]=73;
cos[19421]=73;
cos[19422]=73;
cos[19423]=73;
cos[19424]=73;
cos[19425]=73;
cos[19426]=73;
cos[19427]=73;
cos[19428]=73;
cos[19429]=73;
cos[19430]=73;
cos[19431]=73;
cos[19432]=73;
cos[19433]=73;
cos[19434]=73;
cos[19435]=73;
cos[19436]=73;
cos[19437]=73;
cos[19438]=73;
cos[19439]=73;
cos[19440]=73;
cos[19441]=73;
cos[19442]=73;
cos[19443]=73;
cos[19444]=73;
cos[19445]=73;
cos[19446]=73;
cos[19447]=73;
cos[19448]=73;
cos[19449]=73;
cos[19450]=74;
cos[19451]=74;
cos[19452]=74;
cos[19453]=74;
cos[19454]=74;
cos[19455]=74;
cos[19456]=74;
cos[19457]=74;
cos[19458]=74;
cos[19459]=74;
cos[19460]=74;
cos[19461]=74;
cos[19462]=74;
cos[19463]=74;
cos[19464]=74;
cos[19465]=74;
cos[19466]=74;
cos[19467]=74;
cos[19468]=74;
cos[19469]=74;
cos[19470]=74;
cos[19471]=74;
cos[19472]=74;
cos[19473]=74;
cos[19474]=74;
cos[19475]=74;
cos[19476]=74;
cos[19477]=74;
cos[19478]=74;
cos[19479]=74;
cos[19480]=74;
cos[19481]=74;
cos[19482]=74;
cos[19483]=74;
cos[19484]=74;
cos[19485]=74;
cos[19486]=74;
cos[19487]=74;
cos[19488]=74;
cos[19489]=74;
cos[19490]=74;
cos[19491]=74;
cos[19492]=74;
cos[19493]=74;
cos[19494]=74;
cos[19495]=74;
cos[19496]=74;
cos[19497]=74;
cos[19498]=74;
cos[19499]=74;
cos[19500]=74;
cos[19501]=74;
cos[19502]=74;
cos[19503]=74;
cos[19504]=74;
cos[19505]=74;
cos[19506]=74;
cos[19507]=74;
cos[19508]=74;
cos[19509]=74;
cos[19510]=74;
cos[19511]=74;
cos[19512]=74;
cos[19513]=74;
cos[19514]=75;
cos[19515]=75;
cos[19516]=75;
cos[19517]=75;
cos[19518]=75;
cos[19519]=75;
cos[19520]=75;
cos[19521]=75;
cos[19522]=75;
cos[19523]=75;
cos[19524]=75;
cos[19525]=75;
cos[19526]=75;
cos[19527]=75;
cos[19528]=75;
cos[19529]=75;
cos[19530]=75;
cos[19531]=75;
cos[19532]=75;
cos[19533]=75;
cos[19534]=75;
cos[19535]=75;
cos[19536]=75;
cos[19537]=75;
cos[19538]=75;
cos[19539]=75;
cos[19540]=75;
cos[19541]=75;
cos[19542]=75;
cos[19543]=75;
cos[19544]=75;
cos[19545]=75;
cos[19546]=75;
cos[19547]=75;
cos[19548]=75;
cos[19549]=75;
cos[19550]=75;
cos[19551]=75;
cos[19552]=75;
cos[19553]=75;
cos[19554]=75;
cos[19555]=75;
cos[19556]=75;
cos[19557]=75;
cos[19558]=75;
cos[19559]=75;
cos[19560]=75;
cos[19561]=75;
cos[19562]=75;
cos[19563]=75;
cos[19564]=75;
cos[19565]=75;
cos[19566]=75;
cos[19567]=75;
cos[19568]=75;
cos[19569]=75;
cos[19570]=75;
cos[19571]=75;
cos[19572]=75;
cos[19573]=75;
cos[19574]=75;
cos[19575]=75;
cos[19576]=75;
cos[19577]=75;
cos[19578]=75;
cos[19579]=75;
cos[19580]=75;
cos[19581]=75;
cos[19582]=75;
cos[19583]=75;
cos[19584]=75;
cos[19585]=75;
cos[19586]=75;
cos[19587]=76;
cos[19588]=76;
cos[19589]=76;
cos[19590]=76;
cos[19591]=76;
cos[19592]=76;
cos[19593]=76;
cos[19594]=76;
cos[19595]=76;
cos[19596]=76;
cos[19597]=76;
cos[19598]=76;
cos[19599]=76;
cos[19600]=76;
cos[19601]=76;
cos[19602]=76;
cos[19603]=76;
cos[19604]=76;
cos[19605]=76;
cos[19606]=76;
cos[19607]=76;
cos[19608]=76;
cos[19609]=76;
cos[19610]=76;
cos[19611]=76;
cos[19612]=76;
cos[19613]=76;
cos[19614]=76;
cos[19615]=76;
cos[19616]=76;
cos[19617]=76;
cos[19618]=76;
cos[19619]=76;
cos[19620]=76;
cos[19621]=76;
cos[19622]=76;
cos[19623]=76;
cos[19624]=76;
cos[19625]=76;
cos[19626]=76;
cos[19627]=76;
cos[19628]=76;
cos[19629]=76;
cos[19630]=76;
cos[19631]=76;
cos[19632]=76;
cos[19633]=76;
cos[19634]=76;
cos[19635]=76;
cos[19636]=76;
cos[19637]=76;
cos[19638]=76;
cos[19639]=76;
cos[19640]=76;
cos[19641]=76;
cos[19642]=76;
cos[19643]=76;
cos[19644]=76;
cos[19645]=76;
cos[19646]=76;
cos[19647]=76;
cos[19648]=76;
cos[19649]=76;
cos[19650]=76;
cos[19651]=76;
cos[19652]=76;
cos[19653]=76;
cos[19654]=76;
cos[19655]=76;
cos[19656]=76;
cos[19657]=76;
cos[19658]=76;
cos[19659]=76;
cos[19660]=76;
cos[19661]=76;
cos[19662]=76;
cos[19663]=76;
cos[19664]=76;
cos[19665]=76;
cos[19666]=76;
cos[19667]=76;
cos[19668]=76;
cos[19669]=76;
cos[19670]=76;
cos[19671]=76;
cos[19672]=76;
cos[19673]=76;
cos[19674]=76;
cos[19675]=77;
cos[19676]=77;
cos[19677]=77;
cos[19678]=77;
cos[19679]=77;
cos[19680]=77;
cos[19681]=77;
cos[19682]=77;
cos[19683]=77;
cos[19684]=77;
cos[19685]=77;
cos[19686]=77;
cos[19687]=77;
cos[19688]=77;
cos[19689]=77;
cos[19690]=77;
cos[19691]=77;
cos[19692]=77;
cos[19693]=77;
cos[19694]=77;
cos[19695]=77;
cos[19696]=77;
cos[19697]=77;
cos[19698]=77;
cos[19699]=77;
cos[19700]=77;
cos[19701]=77;
cos[19702]=77;
cos[19703]=77;
cos[19704]=77;
cos[19705]=77;
cos[19706]=77;
cos[19707]=77;
cos[19708]=77;
cos[19709]=77;
cos[19710]=77;
cos[19711]=77;
cos[19712]=77;
cos[19713]=77;
cos[19714]=77;
cos[19715]=77;
cos[19716]=77;
cos[19717]=77;
cos[19718]=77;
cos[19719]=77;
cos[19720]=77;
cos[19721]=77;
cos[19722]=77;
cos[19723]=77;
cos[19724]=77;
cos[19725]=77;
cos[19726]=77;
cos[19727]=77;
cos[19728]=77;
cos[19729]=77;
cos[19730]=77;
cos[19731]=77;
cos[19732]=77;
cos[19733]=77;
cos[19734]=77;
cos[19735]=77;
cos[19736]=77;
cos[19737]=77;
cos[19738]=77;
cos[19739]=77;
cos[19740]=77;
cos[19741]=77;
cos[19742]=77;
cos[19743]=77;
cos[19744]=77;
cos[19745]=77;
cos[19746]=77;
cos[19747]=77;
cos[19748]=77;
cos[19749]=77;
cos[19750]=77;
cos[19751]=77;
cos[19752]=77;
cos[19753]=77;
cos[19754]=77;
cos[19755]=77;
cos[19756]=77;
cos[19757]=77;
cos[19758]=77;
cos[19759]=77;
cos[19760]=77;
cos[19761]=77;
cos[19762]=77;
cos[19763]=77;
cos[19764]=77;
cos[19765]=77;
cos[19766]=77;
cos[19767]=77;
cos[19768]=77;
cos[19769]=77;
cos[19770]=77;
cos[19771]=77;
cos[19772]=77;
cos[19773]=77;
cos[19774]=77;
cos[19775]=77;
cos[19776]=77;
cos[19777]=77;
cos[19778]=77;
cos[19779]=77;
cos[19780]=77;
cos[19781]=77;
cos[19782]=77;
cos[19783]=77;
cos[19784]=77;
cos[19785]=77;
cos[19786]=77;
cos[19787]=77;
cos[19788]=77;
cos[19789]=77;
cos[19790]=77;
cos[19791]=77;
cos[19792]=77;
cos[19793]=77;
cos[19794]=77;
cos[19795]=77;
cos[19796]=77;
cos[19797]=77;
cos[19798]=77;
cos[19799]=78;
cos[19800]=78;
cos[19801]=78;
cos[19802]=78;
cos[19803]=78;
cos[19804]=78;
cos[19805]=78;
cos[19806]=78;
cos[19807]=78;
cos[19808]=78;
cos[19809]=78;
cos[19810]=78;
cos[19811]=78;
cos[19812]=78;
cos[19813]=78;
cos[19814]=78;
cos[19815]=78;
cos[19816]=78;
cos[19817]=78;
cos[19818]=78;
cos[19819]=78;
cos[19820]=78;
cos[19821]=78;
cos[19822]=78;
cos[19823]=78;
cos[19824]=78;
cos[19825]=78;
cos[19826]=78;
cos[19827]=78;
cos[19828]=78;
cos[19829]=78;
cos[19830]=78;
cos[19831]=78;
cos[19832]=78;
cos[19833]=78;
cos[19834]=78;
cos[19835]=78;
cos[19836]=78;
cos[19837]=78;
cos[19838]=78;
cos[19839]=78;
cos[19840]=78;
cos[19841]=78;
cos[19842]=78;
cos[19843]=78;
cos[19844]=78;
cos[19845]=78;
cos[19846]=78;
cos[19847]=78;
cos[19848]=78;
cos[19849]=78;
cos[19850]=78;
cos[19851]=78;
cos[19852]=78;
cos[19853]=78;
cos[19854]=78;
cos[19855]=78;
cos[19856]=78;
cos[19857]=78;
cos[19858]=78;
cos[19859]=78;
cos[19860]=78;
cos[19861]=78;
cos[19862]=78;
cos[19863]=78;
cos[19864]=78;
cos[19865]=78;
cos[19866]=78;
cos[19867]=78;
cos[19868]=78;
cos[19869]=78;
cos[19870]=78;
cos[19871]=78;
cos[19872]=78;
cos[19873]=78;
cos[19874]=78;
cos[19875]=78;
cos[19876]=78;
cos[19877]=78;
cos[19878]=78;
cos[19879]=78;
cos[19880]=78;
cos[19881]=78;
cos[19882]=78;
cos[19883]=78;
cos[19884]=78;
cos[19885]=78;
cos[19886]=78;
cos[19887]=78;
cos[19888]=78;
cos[19889]=78;
cos[19890]=78;
cos[19891]=78;
cos[19892]=78;
cos[19893]=78;
cos[19894]=78;
cos[19895]=78;
cos[19896]=78;
cos[19897]=78;
cos[19898]=78;
cos[19899]=78;
cos[19900]=78;
cos[19901]=78;
cos[19902]=78;
cos[19903]=78;
cos[19904]=78;
cos[19905]=78;
cos[19906]=78;
cos[19907]=78;
cos[19908]=78;
cos[19909]=78;
cos[19910]=78;
cos[19911]=78;
cos[19912]=78;
cos[19913]=78;
cos[19914]=78;
cos[19915]=78;
cos[19916]=78;
cos[19917]=78;
cos[19918]=78;
cos[19919]=78;
cos[19920]=78;
cos[19921]=78;
cos[19922]=78;
cos[19923]=78;
cos[19924]=78;
cos[19925]=78;
cos[19926]=78;
cos[19927]=78;
cos[19928]=78;
cos[19929]=78;
cos[19930]=78;
cos[19931]=78;
cos[19932]=78;
cos[19933]=78;
cos[19934]=78;
cos[19935]=78;
cos[19936]=78;
cos[19937]=78;
cos[19938]=78;
cos[19939]=78;
cos[19940]=78;
cos[19941]=78;
cos[19942]=78;
cos[19943]=78;
cos[19944]=78;
cos[19945]=78;
cos[19946]=78;
cos[19947]=78;
cos[19948]=78;
cos[19949]=78;
cos[19950]=78;
cos[19951]=78;
cos[19952]=78;
cos[19953]=78;
cos[19954]=78;
cos[19955]=78;
cos[19956]=78;
cos[19957]=78;
cos[19958]=78;
cos[19959]=78;
cos[19960]=78;
cos[19961]=78;
cos[19962]=78;
cos[19963]=78;
cos[19964]=78;
cos[19965]=78;
cos[19966]=78;
cos[19967]=78;
cos[19968]=78;
cos[19969]=78;
cos[19970]=78;
cos[19971]=78;
cos[19972]=78;
cos[19973]=78;
cos[19974]=78;
cos[19975]=78;
cos[19976]=78;
cos[19977]=78;
cos[19978]=78;
cos[19979]=78;
cos[19980]=78;
cos[19981]=78;
cos[19982]=78;
cos[19983]=78;
cos[19984]=78;
cos[19985]=78;
cos[19986]=78;
cos[19987]=78;
cos[19988]=78;
cos[19989]=78;
cos[19990]=78;
cos[19991]=78;
cos[19992]=78;
cos[19993]=78;
cos[19994]=78;
cos[19995]=78;
cos[19996]=78;
cos[19997]=78;
cos[19998]=78;
cos[19999]=78;
cos[20000]=78;
cos[20001]=78;
cos[20002]=78;
cos[20003]=78;
cos[20004]=78;
cos[20005]=78;
cos[20006]=78;
cos[20007]=78;
cos[20008]=78;
cos[20009]=78;
cos[20010]=78;
cos[20011]=78;
cos[20012]=78;
cos[20013]=78;
cos[20014]=78;
cos[20015]=78;
cos[20016]=78;
cos[20017]=78;
cos[20018]=78;
cos[20019]=78;
cos[20020]=78;
cos[20021]=78;
cos[20022]=78;
cos[20023]=78;
cos[20024]=78;
cos[20025]=78;
cos[20026]=78;
cos[20027]=78;
cos[20028]=78;
cos[20029]=78;
cos[20030]=78;
cos[20031]=78;
cos[20032]=78;
cos[20033]=78;
cos[20034]=78;
cos[20035]=78;
cos[20036]=78;
cos[20037]=78;
cos[20038]=78;
cos[20039]=78;
cos[20040]=78;
cos[20041]=78;
cos[20042]=78;
cos[20043]=78;
cos[20044]=78;
cos[20045]=78;
cos[20046]=78;
cos[20047]=78;
cos[20048]=78;
cos[20049]=78;
cos[20050]=78;
cos[20051]=78;
cos[20052]=78;
cos[20053]=78;
cos[20054]=78;
cos[20055]=78;
cos[20056]=78;
cos[20057]=78;
cos[20058]=78;
cos[20059]=78;
cos[20060]=78;
cos[20061]=78;
cos[20062]=78;
cos[20063]=78;
cos[20064]=78;
cos[20065]=78;
cos[20066]=78;
cos[20067]=78;
cos[20068]=78;
cos[20069]=78;
cos[20070]=78;
cos[20071]=78;
cos[20072]=78;
cos[20073]=78;
cos[20074]=78;
cos[20075]=78;
cos[20076]=78;
cos[20077]=78;
cos[20078]=78;
cos[20079]=78;
cos[20080]=78;
cos[20081]=78;
cos[20082]=78;
cos[20083]=78;
cos[20084]=78;
cos[20085]=78;
cos[20086]=78;
cos[20087]=78;
cos[20088]=78;
cos[20089]=78;
cos[20090]=78;
cos[20091]=78;
cos[20092]=78;
cos[20093]=78;
cos[20094]=78;
cos[20095]=78;
cos[20096]=78;
cos[20097]=78;
cos[20098]=78;
cos[20099]=78;
cos[20100]=78;
cos[20101]=78;
cos[20102]=78;
cos[20103]=78;
cos[20104]=78;
cos[20105]=78;
cos[20106]=78;
cos[20107]=78;
cos[20108]=78;
cos[20109]=78;
cos[20110]=78;
cos[20111]=78;
cos[20112]=78;
cos[20113]=78;
cos[20114]=78;
cos[20115]=78;
cos[20116]=78;
cos[20117]=78;
cos[20118]=78;
cos[20119]=78;
cos[20120]=78;
cos[20121]=78;
cos[20122]=78;
cos[20123]=78;
cos[20124]=78;
cos[20125]=78;
cos[20126]=78;
cos[20127]=78;
cos[20128]=78;
cos[20129]=78;
cos[20130]=78;
cos[20131]=78;
cos[20132]=78;
cos[20133]=78;
cos[20134]=78;
cos[20135]=78;
cos[20136]=78;
cos[20137]=78;
cos[20138]=78;
cos[20139]=78;
cos[20140]=78;
cos[20141]=78;
cos[20142]=78;
cos[20143]=78;
cos[20144]=78;
cos[20145]=78;
cos[20146]=78;
cos[20147]=78;
cos[20148]=78;
cos[20149]=78;
cos[20150]=78;
cos[20151]=78;
cos[20152]=78;
cos[20153]=78;
cos[20154]=78;
cos[20155]=78;
cos[20156]=78;
cos[20157]=78;
cos[20158]=78;
cos[20159]=78;
cos[20160]=78;
cos[20161]=78;
cos[20162]=78;
cos[20163]=78;
cos[20164]=78;
cos[20165]=78;
cos[20166]=78;
cos[20167]=78;
cos[20168]=78;
cos[20169]=78;
cos[20170]=78;
cos[20171]=78;
cos[20172]=78;
cos[20173]=78;
cos[20174]=78;
cos[20175]=78;
cos[20176]=78;
cos[20177]=78;
cos[20178]=78;
cos[20179]=78;
cos[20180]=78;
cos[20181]=78;
cos[20182]=78;
cos[20183]=78;
cos[20184]=78;
cos[20185]=78;
cos[20186]=78;
cos[20187]=78;
cos[20188]=78;
cos[20189]=78;
cos[20190]=78;
cos[20191]=78;
cos[20192]=78;
cos[20193]=78;
cos[20194]=78;
cos[20195]=78;
cos[20196]=78;
cos[20197]=78;
cos[20198]=78;
cos[20199]=78;
cos[20200]=78;
cos[20201]=78;
cos[20202]=77;
cos[20203]=77;
cos[20204]=77;
cos[20205]=77;
cos[20206]=77;
cos[20207]=77;
cos[20208]=77;
cos[20209]=77;
cos[20210]=77;
cos[20211]=77;
cos[20212]=77;
cos[20213]=77;
cos[20214]=77;
cos[20215]=77;
cos[20216]=77;
cos[20217]=77;
cos[20218]=77;
cos[20219]=77;
cos[20220]=77;
cos[20221]=77;
cos[20222]=77;
cos[20223]=77;
cos[20224]=77;
cos[20225]=77;
cos[20226]=77;
cos[20227]=77;
cos[20228]=77;
cos[20229]=77;
cos[20230]=77;
cos[20231]=77;
cos[20232]=77;
cos[20233]=77;
cos[20234]=77;
cos[20235]=77;
cos[20236]=77;
cos[20237]=77;
cos[20238]=77;
cos[20239]=77;
cos[20240]=77;
cos[20241]=77;
cos[20242]=77;
cos[20243]=77;
cos[20244]=77;
cos[20245]=77;
cos[20246]=77;
cos[20247]=77;
cos[20248]=77;
cos[20249]=77;
cos[20250]=77;
cos[20251]=77;
cos[20252]=77;
cos[20253]=77;
cos[20254]=77;
cos[20255]=77;
cos[20256]=77;
cos[20257]=77;
cos[20258]=77;
cos[20259]=77;
cos[20260]=77;
cos[20261]=77;
cos[20262]=77;
cos[20263]=77;
cos[20264]=77;
cos[20265]=77;
cos[20266]=77;
cos[20267]=77;
cos[20268]=77;
cos[20269]=77;
cos[20270]=77;
cos[20271]=77;
cos[20272]=77;
cos[20273]=77;
cos[20274]=77;
cos[20275]=77;
cos[20276]=77;
cos[20277]=77;
cos[20278]=77;
cos[20279]=77;
cos[20280]=77;
cos[20281]=77;
cos[20282]=77;
cos[20283]=77;
cos[20284]=77;
cos[20285]=77;
cos[20286]=77;
cos[20287]=77;
cos[20288]=77;
cos[20289]=77;
cos[20290]=77;
cos[20291]=77;
cos[20292]=77;
cos[20293]=77;
cos[20294]=77;
cos[20295]=77;
cos[20296]=77;
cos[20297]=77;
cos[20298]=77;
cos[20299]=77;
cos[20300]=77;
cos[20301]=77;
cos[20302]=77;
cos[20303]=77;
cos[20304]=77;
cos[20305]=77;
cos[20306]=77;
cos[20307]=77;
cos[20308]=77;
cos[20309]=77;
cos[20310]=77;
cos[20311]=77;
cos[20312]=77;
cos[20313]=77;
cos[20314]=77;
cos[20315]=77;
cos[20316]=77;
cos[20317]=77;
cos[20318]=77;
cos[20319]=77;
cos[20320]=77;
cos[20321]=77;
cos[20322]=77;
cos[20323]=77;
cos[20324]=77;
cos[20325]=77;
cos[20326]=76;
cos[20327]=76;
cos[20328]=76;
cos[20329]=76;
cos[20330]=76;
cos[20331]=76;
cos[20332]=76;
cos[20333]=76;
cos[20334]=76;
cos[20335]=76;
cos[20336]=76;
cos[20337]=76;
cos[20338]=76;
cos[20339]=76;
cos[20340]=76;
cos[20341]=76;
cos[20342]=76;
cos[20343]=76;
cos[20344]=76;
cos[20345]=76;
cos[20346]=76;
cos[20347]=76;
cos[20348]=76;
cos[20349]=76;
cos[20350]=76;
cos[20351]=76;
cos[20352]=76;
cos[20353]=76;
cos[20354]=76;
cos[20355]=76;
cos[20356]=76;
cos[20357]=76;
cos[20358]=76;
cos[20359]=76;
cos[20360]=76;
cos[20361]=76;
cos[20362]=76;
cos[20363]=76;
cos[20364]=76;
cos[20365]=76;
cos[20366]=76;
cos[20367]=76;
cos[20368]=76;
cos[20369]=76;
cos[20370]=76;
cos[20371]=76;
cos[20372]=76;
cos[20373]=76;
cos[20374]=76;
cos[20375]=76;
cos[20376]=76;
cos[20377]=76;
cos[20378]=76;
cos[20379]=76;
cos[20380]=76;
cos[20381]=76;
cos[20382]=76;
cos[20383]=76;
cos[20384]=76;
cos[20385]=76;
cos[20386]=76;
cos[20387]=76;
cos[20388]=76;
cos[20389]=76;
cos[20390]=76;
cos[20391]=76;
cos[20392]=76;
cos[20393]=76;
cos[20394]=76;
cos[20395]=76;
cos[20396]=76;
cos[20397]=76;
cos[20398]=76;
cos[20399]=76;
cos[20400]=76;
cos[20401]=76;
cos[20402]=76;
cos[20403]=76;
cos[20404]=76;
cos[20405]=76;
cos[20406]=76;
cos[20407]=76;
cos[20408]=76;
cos[20409]=76;
cos[20410]=76;
cos[20411]=76;
cos[20412]=76;
cos[20413]=76;
cos[20414]=75;
cos[20415]=75;
cos[20416]=75;
cos[20417]=75;
cos[20418]=75;
cos[20419]=75;
cos[20420]=75;
cos[20421]=75;
cos[20422]=75;
cos[20423]=75;
cos[20424]=75;
cos[20425]=75;
cos[20426]=75;
cos[20427]=75;
cos[20428]=75;
cos[20429]=75;
cos[20430]=75;
cos[20431]=75;
cos[20432]=75;
cos[20433]=75;
cos[20434]=75;
cos[20435]=75;
cos[20436]=75;
cos[20437]=75;
cos[20438]=75;
cos[20439]=75;
cos[20440]=75;
cos[20441]=75;
cos[20442]=75;
cos[20443]=75;
cos[20444]=75;
cos[20445]=75;
cos[20446]=75;
cos[20447]=75;
cos[20448]=75;
cos[20449]=75;
cos[20450]=75;
cos[20451]=75;
cos[20452]=75;
cos[20453]=75;
cos[20454]=75;
cos[20455]=75;
cos[20456]=75;
cos[20457]=75;
cos[20458]=75;
cos[20459]=75;
cos[20460]=75;
cos[20461]=75;
cos[20462]=75;
cos[20463]=75;
cos[20464]=75;
cos[20465]=75;
cos[20466]=75;
cos[20467]=75;
cos[20468]=75;
cos[20469]=75;
cos[20470]=75;
cos[20471]=75;
cos[20472]=75;
cos[20473]=75;
cos[20474]=75;
cos[20475]=75;
cos[20476]=75;
cos[20477]=75;
cos[20478]=75;
cos[20479]=75;
cos[20480]=75;
cos[20481]=75;
cos[20482]=75;
cos[20483]=75;
cos[20484]=75;
cos[20485]=75;
cos[20486]=75;
cos[20487]=74;
cos[20488]=74;
cos[20489]=74;
cos[20490]=74;
cos[20491]=74;
cos[20492]=74;
cos[20493]=74;
cos[20494]=74;
cos[20495]=74;
cos[20496]=74;
cos[20497]=74;
cos[20498]=74;
cos[20499]=74;
cos[20500]=74;
cos[20501]=74;
cos[20502]=74;
cos[20503]=74;
cos[20504]=74;
cos[20505]=74;
cos[20506]=74;
cos[20507]=74;
cos[20508]=74;
cos[20509]=74;
cos[20510]=74;
cos[20511]=74;
cos[20512]=74;
cos[20513]=74;
cos[20514]=74;
cos[20515]=74;
cos[20516]=74;
cos[20517]=74;
cos[20518]=74;
cos[20519]=74;
cos[20520]=74;
cos[20521]=74;
cos[20522]=74;
cos[20523]=74;
cos[20524]=74;
cos[20525]=74;
cos[20526]=74;
cos[20527]=74;
cos[20528]=74;
cos[20529]=74;
cos[20530]=74;
cos[20531]=74;
cos[20532]=74;
cos[20533]=74;
cos[20534]=74;
cos[20535]=74;
cos[20536]=74;
cos[20537]=74;
cos[20538]=74;
cos[20539]=74;
cos[20540]=74;
cos[20541]=74;
cos[20542]=74;
cos[20543]=74;
cos[20544]=74;
cos[20545]=74;
cos[20546]=74;
cos[20547]=74;
cos[20548]=74;
cos[20549]=74;
cos[20550]=74;
cos[20551]=73;
cos[20552]=73;
cos[20553]=73;
cos[20554]=73;
cos[20555]=73;
cos[20556]=73;
cos[20557]=73;
cos[20558]=73;
cos[20559]=73;
cos[20560]=73;
cos[20561]=73;
cos[20562]=73;
cos[20563]=73;
cos[20564]=73;
cos[20565]=73;
cos[20566]=73;
cos[20567]=73;
cos[20568]=73;
cos[20569]=73;
cos[20570]=73;
cos[20571]=73;
cos[20572]=73;
cos[20573]=73;
cos[20574]=73;
cos[20575]=73;
cos[20576]=73;
cos[20577]=73;
cos[20578]=73;
cos[20579]=73;
cos[20580]=73;
cos[20581]=73;
cos[20582]=73;
cos[20583]=73;
cos[20584]=73;
cos[20585]=73;
cos[20586]=73;
cos[20587]=73;
cos[20588]=73;
cos[20589]=73;
cos[20590]=73;
cos[20591]=73;
cos[20592]=73;
cos[20593]=73;
cos[20594]=73;
cos[20595]=73;
cos[20596]=73;
cos[20597]=73;
cos[20598]=73;
cos[20599]=73;
cos[20600]=73;
cos[20601]=73;
cos[20602]=73;
cos[20603]=73;
cos[20604]=73;
cos[20605]=73;
cos[20606]=73;
cos[20607]=73;
cos[20608]=72;
cos[20609]=72;
cos[20610]=72;
cos[20611]=72;
cos[20612]=72;
cos[20613]=72;
cos[20614]=72;
cos[20615]=72;
cos[20616]=72;
cos[20617]=72;
cos[20618]=72;
cos[20619]=72;
cos[20620]=72;
cos[20621]=72;
cos[20622]=72;
cos[20623]=72;
cos[20624]=72;
cos[20625]=72;
cos[20626]=72;
cos[20627]=72;
cos[20628]=72;
cos[20629]=72;
cos[20630]=72;
cos[20631]=72;
cos[20632]=72;
cos[20633]=72;
cos[20634]=72;
cos[20635]=72;
cos[20636]=72;
cos[20637]=72;
cos[20638]=72;
cos[20639]=72;
cos[20640]=72;
cos[20641]=72;
cos[20642]=72;
cos[20643]=72;
cos[20644]=72;
cos[20645]=72;
cos[20646]=72;
cos[20647]=72;
cos[20648]=72;
cos[20649]=72;
cos[20650]=72;
cos[20651]=72;
cos[20652]=72;
cos[20653]=72;
cos[20654]=72;
cos[20655]=72;
cos[20656]=72;
cos[20657]=72;
cos[20658]=72;
cos[20659]=72;
cos[20660]=72;
cos[20661]=71;
cos[20662]=71;
cos[20663]=71;
cos[20664]=71;
cos[20665]=71;
cos[20666]=71;
cos[20667]=71;
cos[20668]=71;
cos[20669]=71;
cos[20670]=71;
cos[20671]=71;
cos[20672]=71;
cos[20673]=71;
cos[20674]=71;
cos[20675]=71;
cos[20676]=71;
cos[20677]=71;
cos[20678]=71;
cos[20679]=71;
cos[20680]=71;
cos[20681]=71;
cos[20682]=71;
cos[20683]=71;
cos[20684]=71;
cos[20685]=71;
cos[20686]=71;
cos[20687]=71;
cos[20688]=71;
cos[20689]=71;
cos[20690]=71;
cos[20691]=71;
cos[20692]=71;
cos[20693]=71;
cos[20694]=71;
cos[20695]=71;
cos[20696]=71;
cos[20697]=71;
cos[20698]=71;
cos[20699]=71;
cos[20700]=71;
cos[20701]=71;
cos[20702]=71;
cos[20703]=71;
cos[20704]=71;
cos[20705]=71;
cos[20706]=71;
cos[20707]=71;
cos[20708]=71;
cos[20709]=71;
cos[20710]=70;
cos[20711]=70;
cos[20712]=70;
cos[20713]=70;
cos[20714]=70;
cos[20715]=70;
cos[20716]=70;
cos[20717]=70;
cos[20718]=70;
cos[20719]=70;
cos[20720]=70;
cos[20721]=70;
cos[20722]=70;
cos[20723]=70;
cos[20724]=70;
cos[20725]=70;
cos[20726]=70;
cos[20727]=70;
cos[20728]=70;
cos[20729]=70;
cos[20730]=70;
cos[20731]=70;
cos[20732]=70;
cos[20733]=70;
cos[20734]=70;
cos[20735]=70;
cos[20736]=70;
cos[20737]=70;
cos[20738]=70;
cos[20739]=70;
cos[20740]=70;
cos[20741]=70;
cos[20742]=70;
cos[20743]=70;
cos[20744]=70;
cos[20745]=70;
cos[20746]=70;
cos[20747]=70;
cos[20748]=70;
cos[20749]=70;
cos[20750]=70;
cos[20751]=70;
cos[20752]=70;
cos[20753]=70;
cos[20754]=70;
cos[20755]=69;
cos[20756]=69;
cos[20757]=69;
cos[20758]=69;
cos[20759]=69;
cos[20760]=69;
cos[20761]=69;
cos[20762]=69;
cos[20763]=69;
cos[20764]=69;
cos[20765]=69;
cos[20766]=69;
cos[20767]=69;
cos[20768]=69;
cos[20769]=69;
cos[20770]=69;
cos[20771]=69;
cos[20772]=69;
cos[20773]=69;
cos[20774]=69;
cos[20775]=69;
cos[20776]=69;
cos[20777]=69;
cos[20778]=69;
cos[20779]=69;
cos[20780]=69;
cos[20781]=69;
cos[20782]=69;
cos[20783]=69;
cos[20784]=69;
cos[20785]=69;
cos[20786]=69;
cos[20787]=69;
cos[20788]=69;
cos[20789]=69;
cos[20790]=69;
cos[20791]=69;
cos[20792]=69;
cos[20793]=69;
cos[20794]=69;
cos[20795]=69;
cos[20796]=69;
cos[20797]=69;
cos[20798]=69;
cos[20799]=68;
cos[20800]=68;
cos[20801]=68;
cos[20802]=68;
cos[20803]=68;
cos[20804]=68;
cos[20805]=68;
cos[20806]=68;
cos[20807]=68;
cos[20808]=68;
cos[20809]=68;
cos[20810]=68;
cos[20811]=68;
cos[20812]=68;
cos[20813]=68;
cos[20814]=68;
cos[20815]=68;
cos[20816]=68;
cos[20817]=68;
cos[20818]=68;
cos[20819]=68;
cos[20820]=68;
cos[20821]=68;
cos[20822]=68;
cos[20823]=68;
cos[20824]=68;
cos[20825]=68;
cos[20826]=68;
cos[20827]=68;
cos[20828]=68;
cos[20829]=68;
cos[20830]=68;
cos[20831]=68;
cos[20832]=68;
cos[20833]=68;
cos[20834]=68;
cos[20835]=68;
cos[20836]=68;
cos[20837]=68;
cos[20838]=68;
cos[20839]=68;
cos[20840]=67;
cos[20841]=67;
cos[20842]=67;
cos[20843]=67;
cos[20844]=67;
cos[20845]=67;
cos[20846]=67;
cos[20847]=67;
cos[20848]=67;
cos[20849]=67;
cos[20850]=67;
cos[20851]=67;
cos[20852]=67;
cos[20853]=67;
cos[20854]=67;
cos[20855]=67;
cos[20856]=67;
cos[20857]=67;
cos[20858]=67;
cos[20859]=67;
cos[20860]=67;
cos[20861]=67;
cos[20862]=67;
cos[20863]=67;
cos[20864]=67;
cos[20865]=67;
cos[20866]=67;
cos[20867]=67;
cos[20868]=67;
cos[20869]=67;
cos[20870]=67;
cos[20871]=67;
cos[20872]=67;
cos[20873]=67;
cos[20874]=67;
cos[20875]=67;
cos[20876]=67;
cos[20877]=67;
cos[20878]=67;
cos[20879]=67;
cos[20880]=66;
cos[20881]=66;
cos[20882]=66;
cos[20883]=66;
cos[20884]=66;
cos[20885]=66;
cos[20886]=66;
cos[20887]=66;
cos[20888]=66;
cos[20889]=66;
cos[20890]=66;
cos[20891]=66;
cos[20892]=66;
cos[20893]=66;
cos[20894]=66;
cos[20895]=66;
cos[20896]=66;
cos[20897]=66;
cos[20898]=66;
cos[20899]=66;
cos[20900]=66;
cos[20901]=66;
cos[20902]=66;
cos[20903]=66;
cos[20904]=66;
cos[20905]=66;
cos[20906]=66;
cos[20907]=66;
cos[20908]=66;
cos[20909]=66;
cos[20910]=66;
cos[20911]=66;
cos[20912]=66;
cos[20913]=66;
cos[20914]=66;
cos[20915]=66;
cos[20916]=66;
cos[20917]=66;
cos[20918]=65;
cos[20919]=65;
cos[20920]=65;
cos[20921]=65;
cos[20922]=65;
cos[20923]=65;
cos[20924]=65;
cos[20925]=65;
cos[20926]=65;
cos[20927]=65;
cos[20928]=65;
cos[20929]=65;
cos[20930]=65;
cos[20931]=65;
cos[20932]=65;
cos[20933]=65;
cos[20934]=65;
cos[20935]=65;
cos[20936]=65;
cos[20937]=65;
cos[20938]=65;
cos[20939]=65;
cos[20940]=65;
cos[20941]=65;
cos[20942]=65;
cos[20943]=65;
cos[20944]=65;
cos[20945]=65;
cos[20946]=65;
cos[20947]=65;
cos[20948]=65;
cos[20949]=65;
cos[20950]=65;
cos[20951]=65;
cos[20952]=65;
cos[20953]=65;
cos[20954]=65;
cos[20955]=64;
cos[20956]=64;
cos[20957]=64;
cos[20958]=64;
cos[20959]=64;
cos[20960]=64;
cos[20961]=64;
cos[20962]=64;
cos[20963]=64;
cos[20964]=64;
cos[20965]=64;
cos[20966]=64;
cos[20967]=64;
cos[20968]=64;
cos[20969]=64;
cos[20970]=64;
cos[20971]=64;
cos[20972]=64;
cos[20973]=64;
cos[20974]=64;
cos[20975]=64;
cos[20976]=64;
cos[20977]=64;
cos[20978]=64;
cos[20979]=64;
cos[20980]=64;
cos[20981]=64;
cos[20982]=64;
cos[20983]=64;
cos[20984]=64;
cos[20985]=64;
cos[20986]=64;
cos[20987]=64;
cos[20988]=64;
cos[20989]=64;
cos[20990]=63;
cos[20991]=63;
cos[20992]=63;
cos[20993]=63;
cos[20994]=63;
cos[20995]=63;
cos[20996]=63;
cos[20997]=63;
cos[20998]=63;
cos[20999]=63;
cos[21000]=63;
cos[21001]=63;
cos[21002]=63;
cos[21003]=63;
cos[21004]=63;
cos[21005]=63;
cos[21006]=63;
cos[21007]=63;
cos[21008]=63;
cos[21009]=63;
cos[21010]=63;
cos[21011]=63;
cos[21012]=63;
cos[21013]=63;
cos[21014]=63;
cos[21015]=63;
cos[21016]=63;
cos[21017]=63;
cos[21018]=63;
cos[21019]=63;
cos[21020]=63;
cos[21021]=63;
cos[21022]=63;
cos[21023]=63;
cos[21024]=63;
cos[21025]=62;
cos[21026]=62;
cos[21027]=62;
cos[21028]=62;
cos[21029]=62;
cos[21030]=62;
cos[21031]=62;
cos[21032]=62;
cos[21033]=62;
cos[21034]=62;
cos[21035]=62;
cos[21036]=62;
cos[21037]=62;
cos[21038]=62;
cos[21039]=62;
cos[21040]=62;
cos[21041]=62;
cos[21042]=62;
cos[21043]=62;
cos[21044]=62;
cos[21045]=62;
cos[21046]=62;
cos[21047]=62;
cos[21048]=62;
cos[21049]=62;
cos[21050]=62;
cos[21051]=62;
cos[21052]=62;
cos[21053]=62;
cos[21054]=62;
cos[21055]=62;
cos[21056]=62;
cos[21057]=62;
cos[21058]=61;
cos[21059]=61;
cos[21060]=61;
cos[21061]=61;
cos[21062]=61;
cos[21063]=61;
cos[21064]=61;
cos[21065]=61;
cos[21066]=61;
cos[21067]=61;
cos[21068]=61;
cos[21069]=61;
cos[21070]=61;
cos[21071]=61;
cos[21072]=61;
cos[21073]=61;
cos[21074]=61;
cos[21075]=61;
cos[21076]=61;
cos[21077]=61;
cos[21078]=61;
cos[21079]=61;
cos[21080]=61;
cos[21081]=61;
cos[21082]=61;
cos[21083]=61;
cos[21084]=61;
cos[21085]=61;
cos[21086]=61;
cos[21087]=61;
cos[21088]=61;
cos[21089]=61;
cos[21090]=61;
cos[21091]=60;
cos[21092]=60;
cos[21093]=60;
cos[21094]=60;
cos[21095]=60;
cos[21096]=60;
cos[21097]=60;
cos[21098]=60;
cos[21099]=60;
cos[21100]=60;
cos[21101]=60;
cos[21102]=60;
cos[21103]=60;
cos[21104]=60;
cos[21105]=60;
cos[21106]=60;
cos[21107]=60;
cos[21108]=60;
cos[21109]=60;
cos[21110]=60;
cos[21111]=60;
cos[21112]=60;
cos[21113]=60;
cos[21114]=60;
cos[21115]=60;
cos[21116]=60;
cos[21117]=60;
cos[21118]=60;
cos[21119]=60;
cos[21120]=60;
cos[21121]=60;
cos[21122]=60;
cos[21123]=59;
cos[21124]=59;
cos[21125]=59;
cos[21126]=59;
cos[21127]=59;
cos[21128]=59;
cos[21129]=59;
cos[21130]=59;
cos[21131]=59;
cos[21132]=59;
cos[21133]=59;
cos[21134]=59;
cos[21135]=59;
cos[21136]=59;
cos[21137]=59;
cos[21138]=59;
cos[21139]=59;
cos[21140]=59;
cos[21141]=59;
cos[21142]=59;
cos[21143]=59;
cos[21144]=59;
cos[21145]=59;
cos[21146]=59;
cos[21147]=59;
cos[21148]=59;
cos[21149]=59;
cos[21150]=59;
cos[21151]=59;
cos[21152]=59;
cos[21153]=59;
cos[21154]=58;
cos[21155]=58;
cos[21156]=58;
cos[21157]=58;
cos[21158]=58;
cos[21159]=58;
cos[21160]=58;
cos[21161]=58;
cos[21162]=58;
cos[21163]=58;
cos[21164]=58;
cos[21165]=58;
cos[21166]=58;
cos[21167]=58;
cos[21168]=58;
cos[21169]=58;
cos[21170]=58;
cos[21171]=58;
cos[21172]=58;
cos[21173]=58;
cos[21174]=58;
cos[21175]=58;
cos[21176]=58;
cos[21177]=58;
cos[21178]=58;
cos[21179]=58;
cos[21180]=58;
cos[21181]=58;
cos[21182]=58;
cos[21183]=58;
cos[21184]=57;
cos[21185]=57;
cos[21186]=57;
cos[21187]=57;
cos[21188]=57;
cos[21189]=57;
cos[21190]=57;
cos[21191]=57;
cos[21192]=57;
cos[21193]=57;
cos[21194]=57;
cos[21195]=57;
cos[21196]=57;
cos[21197]=57;
cos[21198]=57;
cos[21199]=57;
cos[21200]=57;
cos[21201]=57;
cos[21202]=57;
cos[21203]=57;
cos[21204]=57;
cos[21205]=57;
cos[21206]=57;
cos[21207]=57;
cos[21208]=57;
cos[21209]=57;
cos[21210]=57;
cos[21211]=57;
cos[21212]=57;
cos[21213]=57;
cos[21214]=56;
cos[21215]=56;
cos[21216]=56;
cos[21217]=56;
cos[21218]=56;
cos[21219]=56;
cos[21220]=56;
cos[21221]=56;
cos[21222]=56;
cos[21223]=56;
cos[21224]=56;
cos[21225]=56;
cos[21226]=56;
cos[21227]=56;
cos[21228]=56;
cos[21229]=56;
cos[21230]=56;
cos[21231]=56;
cos[21232]=56;
cos[21233]=56;
cos[21234]=56;
cos[21235]=56;
cos[21236]=56;
cos[21237]=56;
cos[21238]=56;
cos[21239]=56;
cos[21240]=56;
cos[21241]=56;
cos[21242]=56;
cos[21243]=55;
cos[21244]=55;
cos[21245]=55;
cos[21246]=55;
cos[21247]=55;
cos[21248]=55;
cos[21249]=55;
cos[21250]=55;
cos[21251]=55;
cos[21252]=55;
cos[21253]=55;
cos[21254]=55;
cos[21255]=55;
cos[21256]=55;
cos[21257]=55;
cos[21258]=55;
cos[21259]=55;
cos[21260]=55;
cos[21261]=55;
cos[21262]=55;
cos[21263]=55;
cos[21264]=55;
cos[21265]=55;
cos[21266]=55;
cos[21267]=55;
cos[21268]=55;
cos[21269]=55;
cos[21270]=55;
cos[21271]=55;
cos[21272]=54;
cos[21273]=54;
cos[21274]=54;
cos[21275]=54;
cos[21276]=54;
cos[21277]=54;
cos[21278]=54;
cos[21279]=54;
cos[21280]=54;
cos[21281]=54;
cos[21282]=54;
cos[21283]=54;
cos[21284]=54;
cos[21285]=54;
cos[21286]=54;
cos[21287]=54;
cos[21288]=54;
cos[21289]=54;
cos[21290]=54;
cos[21291]=54;
cos[21292]=54;
cos[21293]=54;
cos[21294]=54;
cos[21295]=54;
cos[21296]=54;
cos[21297]=54;
cos[21298]=54;
cos[21299]=54;
cos[21300]=53;
cos[21301]=53;
cos[21302]=53;
cos[21303]=53;
cos[21304]=53;
cos[21305]=53;
cos[21306]=53;
cos[21307]=53;
cos[21308]=53;
cos[21309]=53;
cos[21310]=53;
cos[21311]=53;
cos[21312]=53;
cos[21313]=53;
cos[21314]=53;
cos[21315]=53;
cos[21316]=53;
cos[21317]=53;
cos[21318]=53;
cos[21319]=53;
cos[21320]=53;
cos[21321]=53;
cos[21322]=53;
cos[21323]=53;
cos[21324]=53;
cos[21325]=53;
cos[21326]=53;
cos[21327]=53;
cos[21328]=52;
cos[21329]=52;
cos[21330]=52;
cos[21331]=52;
cos[21332]=52;
cos[21333]=52;
cos[21334]=52;
cos[21335]=52;
cos[21336]=52;
cos[21337]=52;
cos[21338]=52;
cos[21339]=52;
cos[21340]=52;
cos[21341]=52;
cos[21342]=52;
cos[21343]=52;
cos[21344]=52;
cos[21345]=52;
cos[21346]=52;
cos[21347]=52;
cos[21348]=52;
cos[21349]=52;
cos[21350]=52;
cos[21351]=52;
cos[21352]=52;
cos[21353]=52;
cos[21354]=52;
cos[21355]=51;
cos[21356]=51;
cos[21357]=51;
cos[21358]=51;
cos[21359]=51;
cos[21360]=51;
cos[21361]=51;
cos[21362]=51;
cos[21363]=51;
cos[21364]=51;
cos[21365]=51;
cos[21366]=51;
cos[21367]=51;
cos[21368]=51;
cos[21369]=51;
cos[21370]=51;
cos[21371]=51;
cos[21372]=51;
cos[21373]=51;
cos[21374]=51;
cos[21375]=51;
cos[21376]=51;
cos[21377]=51;
cos[21378]=51;
cos[21379]=51;
cos[21380]=51;
cos[21381]=51;
cos[21382]=50;
cos[21383]=50;
cos[21384]=50;
cos[21385]=50;
cos[21386]=50;
cos[21387]=50;
cos[21388]=50;
cos[21389]=50;
cos[21390]=50;
cos[21391]=50;
cos[21392]=50;
cos[21393]=50;
cos[21394]=50;
cos[21395]=50;
cos[21396]=50;
cos[21397]=50;
cos[21398]=50;
cos[21399]=50;
cos[21400]=50;
cos[21401]=50;
cos[21402]=50;
cos[21403]=50;
cos[21404]=50;
cos[21405]=50;
cos[21406]=50;
cos[21407]=50;
cos[21408]=49;
cos[21409]=49;
cos[21410]=49;
cos[21411]=49;
cos[21412]=49;
cos[21413]=49;
cos[21414]=49;
cos[21415]=49;
cos[21416]=49;
cos[21417]=49;
cos[21418]=49;
cos[21419]=49;
cos[21420]=49;
cos[21421]=49;
cos[21422]=49;
cos[21423]=49;
cos[21424]=49;
cos[21425]=49;
cos[21426]=49;
cos[21427]=49;
cos[21428]=49;
cos[21429]=49;
cos[21430]=49;
cos[21431]=49;
cos[21432]=49;
cos[21433]=49;
cos[21434]=49;
cos[21435]=48;
cos[21436]=48;
cos[21437]=48;
cos[21438]=48;
cos[21439]=48;
cos[21440]=48;
cos[21441]=48;
cos[21442]=48;
cos[21443]=48;
cos[21444]=48;
cos[21445]=48;
cos[21446]=48;
cos[21447]=48;
cos[21448]=48;
cos[21449]=48;
cos[21450]=48;
cos[21451]=48;
cos[21452]=48;
cos[21453]=48;
cos[21454]=48;
cos[21455]=48;
cos[21456]=48;
cos[21457]=48;
cos[21458]=48;
cos[21459]=48;
cos[21460]=47;
cos[21461]=47;
cos[21462]=47;
cos[21463]=47;
cos[21464]=47;
cos[21465]=47;
cos[21466]=47;
cos[21467]=47;
cos[21468]=47;
cos[21469]=47;
cos[21470]=47;
cos[21471]=47;
cos[21472]=47;
cos[21473]=47;
cos[21474]=47;
cos[21475]=47;
cos[21476]=47;
cos[21477]=47;
cos[21478]=47;
cos[21479]=47;
cos[21480]=47;
cos[21481]=47;
cos[21482]=47;
cos[21483]=47;
cos[21484]=47;
cos[21485]=47;
cos[21486]=46;
cos[21487]=46;
cos[21488]=46;
cos[21489]=46;
cos[21490]=46;
cos[21491]=46;
cos[21492]=46;
cos[21493]=46;
cos[21494]=46;
cos[21495]=46;
cos[21496]=46;
cos[21497]=46;
cos[21498]=46;
cos[21499]=46;
cos[21500]=46;
cos[21501]=46;
cos[21502]=46;
cos[21503]=46;
cos[21504]=46;
cos[21505]=46;
cos[21506]=46;
cos[21507]=46;
cos[21508]=46;
cos[21509]=46;
cos[21510]=46;
cos[21511]=45;
cos[21512]=45;
cos[21513]=45;
cos[21514]=45;
cos[21515]=45;
cos[21516]=45;
cos[21517]=45;
cos[21518]=45;
cos[21519]=45;
cos[21520]=45;
cos[21521]=45;
cos[21522]=45;
cos[21523]=45;
cos[21524]=45;
cos[21525]=45;
cos[21526]=45;
cos[21527]=45;
cos[21528]=45;
cos[21529]=45;
cos[21530]=45;
cos[21531]=45;
cos[21532]=45;
cos[21533]=45;
cos[21534]=45;
cos[21535]=45;
cos[21536]=44;
cos[21537]=44;
cos[21538]=44;
cos[21539]=44;
cos[21540]=44;
cos[21541]=44;
cos[21542]=44;
cos[21543]=44;
cos[21544]=44;
cos[21545]=44;
cos[21546]=44;
cos[21547]=44;
cos[21548]=44;
cos[21549]=44;
cos[21550]=44;
cos[21551]=44;
cos[21552]=44;
cos[21553]=44;
cos[21554]=44;
cos[21555]=44;
cos[21556]=44;
cos[21557]=44;
cos[21558]=44;
cos[21559]=44;
cos[21560]=44;
cos[21561]=43;
cos[21562]=43;
cos[21563]=43;
cos[21564]=43;
cos[21565]=43;
cos[21566]=43;
cos[21567]=43;
cos[21568]=43;
cos[21569]=43;
cos[21570]=43;
cos[21571]=43;
cos[21572]=43;
cos[21573]=43;
cos[21574]=43;
cos[21575]=43;
cos[21576]=43;
cos[21577]=43;
cos[21578]=43;
cos[21579]=43;
cos[21580]=43;
cos[21581]=43;
cos[21582]=43;
cos[21583]=43;
cos[21584]=43;
cos[21585]=42;
cos[21586]=42;
cos[21587]=42;
cos[21588]=42;
cos[21589]=42;
cos[21590]=42;
cos[21591]=42;
cos[21592]=42;
cos[21593]=42;
cos[21594]=42;
cos[21595]=42;
cos[21596]=42;
cos[21597]=42;
cos[21598]=42;
cos[21599]=42;
cos[21600]=42;
cos[21601]=42;
cos[21602]=42;
cos[21603]=42;
cos[21604]=42;
cos[21605]=42;
cos[21606]=42;
cos[21607]=42;
cos[21608]=42;
cos[21609]=41;
cos[21610]=41;
cos[21611]=41;
cos[21612]=41;
cos[21613]=41;
cos[21614]=41;
cos[21615]=41;
cos[21616]=41;
cos[21617]=41;
cos[21618]=41;
cos[21619]=41;
cos[21620]=41;
cos[21621]=41;
cos[21622]=41;
cos[21623]=41;
cos[21624]=41;
cos[21625]=41;
cos[21626]=41;
cos[21627]=41;
cos[21628]=41;
cos[21629]=41;
cos[21630]=41;
cos[21631]=41;
cos[21632]=41;
cos[21633]=40;
cos[21634]=40;
cos[21635]=40;
cos[21636]=40;
cos[21637]=40;
cos[21638]=40;
cos[21639]=40;
cos[21640]=40;
cos[21641]=40;
cos[21642]=40;
cos[21643]=40;
cos[21644]=40;
cos[21645]=40;
cos[21646]=40;
cos[21647]=40;
cos[21648]=40;
cos[21649]=40;
cos[21650]=40;
cos[21651]=40;
cos[21652]=40;
cos[21653]=40;
cos[21654]=40;
cos[21655]=40;
cos[21656]=40;
cos[21657]=39;
cos[21658]=39;
cos[21659]=39;
cos[21660]=39;
cos[21661]=39;
cos[21662]=39;
cos[21663]=39;
cos[21664]=39;
cos[21665]=39;
cos[21666]=39;
cos[21667]=39;
cos[21668]=39;
cos[21669]=39;
cos[21670]=39;
cos[21671]=39;
cos[21672]=39;
cos[21673]=39;
cos[21674]=39;
cos[21675]=39;
cos[21676]=39;
cos[21677]=39;
cos[21678]=39;
cos[21679]=39;
cos[21680]=38;
cos[21681]=38;
cos[21682]=38;
cos[21683]=38;
cos[21684]=38;
cos[21685]=38;
cos[21686]=38;
cos[21687]=38;
cos[21688]=38;
cos[21689]=38;
cos[21690]=38;
cos[21691]=38;
cos[21692]=38;
cos[21693]=38;
cos[21694]=38;
cos[21695]=38;
cos[21696]=38;
cos[21697]=38;
cos[21698]=38;
cos[21699]=38;
cos[21700]=38;
cos[21701]=38;
cos[21702]=38;
cos[21703]=38;
cos[21704]=37;
cos[21705]=37;
cos[21706]=37;
cos[21707]=37;
cos[21708]=37;
cos[21709]=37;
cos[21710]=37;
cos[21711]=37;
cos[21712]=37;
cos[21713]=37;
cos[21714]=37;
cos[21715]=37;
cos[21716]=37;
cos[21717]=37;
cos[21718]=37;
cos[21719]=37;
cos[21720]=37;
cos[21721]=37;
cos[21722]=37;
cos[21723]=37;
cos[21724]=37;
cos[21725]=37;
cos[21726]=37;
cos[21727]=36;
cos[21728]=36;
cos[21729]=36;
cos[21730]=36;
cos[21731]=36;
cos[21732]=36;
cos[21733]=36;
cos[21734]=36;
cos[21735]=36;
cos[21736]=36;
cos[21737]=36;
cos[21738]=36;
cos[21739]=36;
cos[21740]=36;
cos[21741]=36;
cos[21742]=36;
cos[21743]=36;
cos[21744]=36;
cos[21745]=36;
cos[21746]=36;
cos[21747]=36;
cos[21748]=36;
cos[21749]=36;
cos[21750]=35;
cos[21751]=35;
cos[21752]=35;
cos[21753]=35;
cos[21754]=35;
cos[21755]=35;
cos[21756]=35;
cos[21757]=35;
cos[21758]=35;
cos[21759]=35;
cos[21760]=35;
cos[21761]=35;
cos[21762]=35;
cos[21763]=35;
cos[21764]=35;
cos[21765]=35;
cos[21766]=35;
cos[21767]=35;
cos[21768]=35;
cos[21769]=35;
cos[21770]=35;
cos[21771]=35;
cos[21772]=35;
cos[21773]=34;
cos[21774]=34;
cos[21775]=34;
cos[21776]=34;
cos[21777]=34;
cos[21778]=34;
cos[21779]=34;
cos[21780]=34;
cos[21781]=34;
cos[21782]=34;
cos[21783]=34;
cos[21784]=34;
cos[21785]=34;
cos[21786]=34;
cos[21787]=34;
cos[21788]=34;
cos[21789]=34;
cos[21790]=34;
cos[21791]=34;
cos[21792]=34;
cos[21793]=34;
cos[21794]=34;
cos[21795]=33;
cos[21796]=33;
cos[21797]=33;
cos[21798]=33;
cos[21799]=33;
cos[21800]=33;
cos[21801]=33;
cos[21802]=33;
cos[21803]=33;
cos[21804]=33;
cos[21805]=33;
cos[21806]=33;
cos[21807]=33;
cos[21808]=33;
cos[21809]=33;
cos[21810]=33;
cos[21811]=33;
cos[21812]=33;
cos[21813]=33;
cos[21814]=33;
cos[21815]=33;
cos[21816]=33;
cos[21817]=33;
cos[21818]=32;
cos[21819]=32;
cos[21820]=32;
cos[21821]=32;
cos[21822]=32;
cos[21823]=32;
cos[21824]=32;
cos[21825]=32;
cos[21826]=32;
cos[21827]=32;
cos[21828]=32;
cos[21829]=32;
cos[21830]=32;
cos[21831]=32;
cos[21832]=32;
cos[21833]=32;
cos[21834]=32;
cos[21835]=32;
cos[21836]=32;
cos[21837]=32;
cos[21838]=32;
cos[21839]=32;
cos[21840]=31;
cos[21841]=31;
cos[21842]=31;
cos[21843]=31;
cos[21844]=31;
cos[21845]=31;
cos[21846]=31;
cos[21847]=31;
cos[21848]=31;
cos[21849]=31;
cos[21850]=31;
cos[21851]=31;
cos[21852]=31;
cos[21853]=31;
cos[21854]=31;
cos[21855]=31;
cos[21856]=31;
cos[21857]=31;
cos[21858]=31;
cos[21859]=31;
cos[21860]=31;
cos[21861]=31;
cos[21862]=30;
cos[21863]=30;
cos[21864]=30;
cos[21865]=30;
cos[21866]=30;
cos[21867]=30;
cos[21868]=30;
cos[21869]=30;
cos[21870]=30;
cos[21871]=30;
cos[21872]=30;
cos[21873]=30;
cos[21874]=30;
cos[21875]=30;
cos[21876]=30;
cos[21877]=30;
cos[21878]=30;
cos[21879]=30;
cos[21880]=30;
cos[21881]=30;
cos[21882]=30;
cos[21883]=30;
cos[21884]=29;
cos[21885]=29;
cos[21886]=29;
cos[21887]=29;
cos[21888]=29;
cos[21889]=29;
cos[21890]=29;
cos[21891]=29;
cos[21892]=29;
cos[21893]=29;
cos[21894]=29;
cos[21895]=29;
cos[21896]=29;
cos[21897]=29;
cos[21898]=29;
cos[21899]=29;
cos[21900]=29;
cos[21901]=29;
cos[21902]=29;
cos[21903]=29;
cos[21904]=29;
cos[21905]=29;
cos[21906]=28;
cos[21907]=28;
cos[21908]=28;
cos[21909]=28;
cos[21910]=28;
cos[21911]=28;
cos[21912]=28;
cos[21913]=28;
cos[21914]=28;
cos[21915]=28;
cos[21916]=28;
cos[21917]=28;
cos[21918]=28;
cos[21919]=28;
cos[21920]=28;
cos[21921]=28;
cos[21922]=28;
cos[21923]=28;
cos[21924]=28;
cos[21925]=28;
cos[21926]=28;
cos[21927]=28;
cos[21928]=27;
cos[21929]=27;
cos[21930]=27;
cos[21931]=27;
cos[21932]=27;
cos[21933]=27;
cos[21934]=27;
cos[21935]=27;
cos[21936]=27;
cos[21937]=27;
cos[21938]=27;
cos[21939]=27;
cos[21940]=27;
cos[21941]=27;
cos[21942]=27;
cos[21943]=27;
cos[21944]=27;
cos[21945]=27;
cos[21946]=27;
cos[21947]=27;
cos[21948]=27;
cos[21949]=27;
cos[21950]=26;
cos[21951]=26;
cos[21952]=26;
cos[21953]=26;
cos[21954]=26;
cos[21955]=26;
cos[21956]=26;
cos[21957]=26;
cos[21958]=26;
cos[21959]=26;
cos[21960]=26;
cos[21961]=26;
cos[21962]=26;
cos[21963]=26;
cos[21964]=26;
cos[21965]=26;
cos[21966]=26;
cos[21967]=26;
cos[21968]=26;
cos[21969]=26;
cos[21970]=26;
cos[21971]=25;
cos[21972]=25;
cos[21973]=25;
cos[21974]=25;
cos[21975]=25;
cos[21976]=25;
cos[21977]=25;
cos[21978]=25;
cos[21979]=25;
cos[21980]=25;
cos[21981]=25;
cos[21982]=25;
cos[21983]=25;
cos[21984]=25;
cos[21985]=25;
cos[21986]=25;
cos[21987]=25;
cos[21988]=25;
cos[21989]=25;
cos[21990]=25;
cos[21991]=25;
cos[21992]=25;
cos[21993]=24;
cos[21994]=24;
cos[21995]=24;
cos[21996]=24;
cos[21997]=24;
cos[21998]=24;
cos[21999]=24;
cos[22000]=24;
cos[22001]=24;
cos[22002]=24;
cos[22003]=24;
cos[22004]=24;
cos[22005]=24;
cos[22006]=24;
cos[22007]=24;
cos[22008]=24;
cos[22009]=24;
cos[22010]=24;
cos[22011]=24;
cos[22012]=24;
cos[22013]=24;
cos[22014]=23;
cos[22015]=23;
cos[22016]=23;
cos[22017]=23;
cos[22018]=23;
cos[22019]=23;
cos[22020]=23;
cos[22021]=23;
cos[22022]=23;
cos[22023]=23;
cos[22024]=23;
cos[22025]=23;
cos[22026]=23;
cos[22027]=23;
cos[22028]=23;
cos[22029]=23;
cos[22030]=23;
cos[22031]=23;
cos[22032]=23;
cos[22033]=23;
cos[22034]=23;
cos[22035]=23;
cos[22036]=22;
cos[22037]=22;
cos[22038]=22;
cos[22039]=22;
cos[22040]=22;
cos[22041]=22;
cos[22042]=22;
cos[22043]=22;
cos[22044]=22;
cos[22045]=22;
cos[22046]=22;
cos[22047]=22;
cos[22048]=22;
cos[22049]=22;
cos[22050]=22;
cos[22051]=22;
cos[22052]=22;
cos[22053]=22;
cos[22054]=22;
cos[22055]=22;
cos[22056]=22;
cos[22057]=21;
cos[22058]=21;
cos[22059]=21;
cos[22060]=21;
cos[22061]=21;
cos[22062]=21;
cos[22063]=21;
cos[22064]=21;
cos[22065]=21;
cos[22066]=21;
cos[22067]=21;
cos[22068]=21;
cos[22069]=21;
cos[22070]=21;
cos[22071]=21;
cos[22072]=21;
cos[22073]=21;
cos[22074]=21;
cos[22075]=21;
cos[22076]=21;
cos[22077]=21;
cos[22078]=20;
cos[22079]=20;
cos[22080]=20;
cos[22081]=20;
cos[22082]=20;
cos[22083]=20;
cos[22084]=20;
cos[22085]=20;
cos[22086]=20;
cos[22087]=20;
cos[22088]=20;
cos[22089]=20;
cos[22090]=20;
cos[22091]=20;
cos[22092]=20;
cos[22093]=20;
cos[22094]=20;
cos[22095]=20;
cos[22096]=20;
cos[22097]=20;
cos[22098]=20;
cos[22099]=19;
cos[22100]=19;
cos[22101]=19;
cos[22102]=19;
cos[22103]=19;
cos[22104]=19;
cos[22105]=19;
cos[22106]=19;
cos[22107]=19;
cos[22108]=19;
cos[22109]=19;
cos[22110]=19;
cos[22111]=19;
cos[22112]=19;
cos[22113]=19;
cos[22114]=19;
cos[22115]=19;
cos[22116]=19;
cos[22117]=19;
cos[22118]=19;
cos[22119]=19;
cos[22120]=18;
cos[22121]=18;
cos[22122]=18;
cos[22123]=18;
cos[22124]=18;
cos[22125]=18;
cos[22126]=18;
cos[22127]=18;
cos[22128]=18;
cos[22129]=18;
cos[22130]=18;
cos[22131]=18;
cos[22132]=18;
cos[22133]=18;
cos[22134]=18;
cos[22135]=18;
cos[22136]=18;
cos[22137]=18;
cos[22138]=18;
cos[22139]=18;
cos[22140]=18;
cos[22141]=17;
cos[22142]=17;
cos[22143]=17;
cos[22144]=17;
cos[22145]=17;
cos[22146]=17;
cos[22147]=17;
cos[22148]=17;
cos[22149]=17;
cos[22150]=17;
cos[22151]=17;
cos[22152]=17;
cos[22153]=17;
cos[22154]=17;
cos[22155]=17;
cos[22156]=17;
cos[22157]=17;
cos[22158]=17;
cos[22159]=17;
cos[22160]=17;
cos[22161]=17;
cos[22162]=16;
cos[22163]=16;
cos[22164]=16;
cos[22165]=16;
cos[22166]=16;
cos[22167]=16;
cos[22168]=16;
cos[22169]=16;
cos[22170]=16;
cos[22171]=16;
cos[22172]=16;
cos[22173]=16;
cos[22174]=16;
cos[22175]=16;
cos[22176]=16;
cos[22177]=16;
cos[22178]=16;
cos[22179]=16;
cos[22180]=16;
cos[22181]=16;
cos[22182]=16;
cos[22183]=15;
cos[22184]=15;
cos[22185]=15;
cos[22186]=15;
cos[22187]=15;
cos[22188]=15;
cos[22189]=15;
cos[22190]=15;
cos[22191]=15;
cos[22192]=15;
cos[22193]=15;
cos[22194]=15;
cos[22195]=15;
cos[22196]=15;
cos[22197]=15;
cos[22198]=15;
cos[22199]=15;
cos[22200]=15;
cos[22201]=15;
cos[22202]=15;
cos[22203]=14;
cos[22204]=14;
cos[22205]=14;
cos[22206]=14;
cos[22207]=14;
cos[22208]=14;
cos[22209]=14;
cos[22210]=14;
cos[22211]=14;
cos[22212]=14;
cos[22213]=14;
cos[22214]=14;
cos[22215]=14;
cos[22216]=14;
cos[22217]=14;
cos[22218]=14;
cos[22219]=14;
cos[22220]=14;
cos[22221]=14;
cos[22222]=14;
cos[22223]=14;
cos[22224]=13;
cos[22225]=13;
cos[22226]=13;
cos[22227]=13;
cos[22228]=13;
cos[22229]=13;
cos[22230]=13;
cos[22231]=13;
cos[22232]=13;
cos[22233]=13;
cos[22234]=13;
cos[22235]=13;
cos[22236]=13;
cos[22237]=13;
cos[22238]=13;
cos[22239]=13;
cos[22240]=13;
cos[22241]=13;
cos[22242]=13;
cos[22243]=13;
cos[22244]=13;
cos[22245]=12;
cos[22246]=12;
cos[22247]=12;
cos[22248]=12;
cos[22249]=12;
cos[22250]=12;
cos[22251]=12;
cos[22252]=12;
cos[22253]=12;
cos[22254]=12;
cos[22255]=12;
cos[22256]=12;
cos[22257]=12;
cos[22258]=12;
cos[22259]=12;
cos[22260]=12;
cos[22261]=12;
cos[22262]=12;
cos[22263]=12;
cos[22264]=12;
cos[22265]=11;
cos[22266]=11;
cos[22267]=11;
cos[22268]=11;
cos[22269]=11;
cos[22270]=11;
cos[22271]=11;
cos[22272]=11;
cos[22273]=11;
cos[22274]=11;
cos[22275]=11;
cos[22276]=11;
cos[22277]=11;
cos[22278]=11;
cos[22279]=11;
cos[22280]=11;
cos[22281]=11;
cos[22282]=11;
cos[22283]=11;
cos[22284]=11;
cos[22285]=11;
cos[22286]=10;
cos[22287]=10;
cos[22288]=10;
cos[22289]=10;
cos[22290]=10;
cos[22291]=10;
cos[22292]=10;
cos[22293]=10;
cos[22294]=10;
cos[22295]=10;
cos[22296]=10;
cos[22297]=10;
cos[22298]=10;
cos[22299]=10;
cos[22300]=10;
cos[22301]=10;
cos[22302]=10;
cos[22303]=10;
cos[22304]=10;
cos[22305]=10;
cos[22306]=9;
cos[22307]=9;
cos[22308]=9;
cos[22309]=9;
cos[22310]=9;
cos[22311]=9;
cos[22312]=9;
cos[22313]=9;
cos[22314]=9;
cos[22315]=9;
cos[22316]=9;
cos[22317]=9;
cos[22318]=9;
cos[22319]=9;
cos[22320]=9;
cos[22321]=9;
cos[22322]=9;
cos[22323]=9;
cos[22324]=9;
cos[22325]=9;
cos[22326]=9;
cos[22327]=8;
cos[22328]=8;
cos[22329]=8;
cos[22330]=8;
cos[22331]=8;
cos[22332]=8;
cos[22333]=8;
cos[22334]=8;
cos[22335]=8;
cos[22336]=8;
cos[22337]=8;
cos[22338]=8;
cos[22339]=8;
cos[22340]=8;
cos[22341]=8;
cos[22342]=8;
cos[22343]=8;
cos[22344]=8;
cos[22345]=8;
cos[22346]=8;
cos[22347]=7;
cos[22348]=7;
cos[22349]=7;
cos[22350]=7;
cos[22351]=7;
cos[22352]=7;
cos[22353]=7;
cos[22354]=7;
cos[22355]=7;
cos[22356]=7;
cos[22357]=7;
cos[22358]=7;
cos[22359]=7;
cos[22360]=7;
cos[22361]=7;
cos[22362]=7;
cos[22363]=7;
cos[22364]=7;
cos[22365]=7;
cos[22366]=7;
cos[22367]=7;
cos[22368]=6;
cos[22369]=6;
cos[22370]=6;
cos[22371]=6;
cos[22372]=6;
cos[22373]=6;
cos[22374]=6;
cos[22375]=6;
cos[22376]=6;
cos[22377]=6;
cos[22378]=6;
cos[22379]=6;
cos[22380]=6;
cos[22381]=6;
cos[22382]=6;
cos[22383]=6;
cos[22384]=6;
cos[22385]=6;
cos[22386]=6;
cos[22387]=6;
cos[22388]=5;
cos[22389]=5;
cos[22390]=5;
cos[22391]=5;
cos[22392]=5;
cos[22393]=5;
cos[22394]=5;
cos[22395]=5;
cos[22396]=5;
cos[22397]=5;
cos[22398]=5;
cos[22399]=5;
cos[22400]=5;
cos[22401]=5;
cos[22402]=5;
cos[22403]=5;
cos[22404]=5;
cos[22405]=5;
cos[22406]=5;
cos[22407]=5;
cos[22408]=5;
cos[22409]=4;
cos[22410]=4;
cos[22411]=4;
cos[22412]=4;
cos[22413]=4;
cos[22414]=4;
cos[22415]=4;
cos[22416]=4;
cos[22417]=4;
cos[22418]=4;
cos[22419]=4;
cos[22420]=4;
cos[22421]=4;
cos[22422]=4;
cos[22423]=4;
cos[22424]=4;
cos[22425]=4;
cos[22426]=4;
cos[22427]=4;
cos[22428]=4;
cos[22429]=3;
cos[22430]=3;
cos[22431]=3;
cos[22432]=3;
cos[22433]=3;
cos[22434]=3;
cos[22435]=3;
cos[22436]=3;
cos[22437]=3;
cos[22438]=3;
cos[22439]=3;
cos[22440]=3;
cos[22441]=3;
cos[22442]=3;
cos[22443]=3;
cos[22444]=3;
cos[22445]=3;
cos[22446]=3;
cos[22447]=3;
cos[22448]=3;
cos[22449]=3;
cos[22450]=2;
cos[22451]=2;
cos[22452]=2;
cos[22453]=2;
cos[22454]=2;
cos[22455]=2;
cos[22456]=2;
cos[22457]=2;
cos[22458]=2;
cos[22459]=2;
cos[22460]=2;
cos[22461]=2;
cos[22462]=2;
cos[22463]=2;
cos[22464]=2;
cos[22465]=2;
cos[22466]=2;
cos[22467]=2;
cos[22468]=2;
cos[22469]=2;
cos[22470]=1;
cos[22471]=1;
cos[22472]=1;
cos[22473]=1;
cos[22474]=1;
cos[22475]=1;
cos[22476]=1;
cos[22477]=1;
cos[22478]=1;
cos[22479]=1;
cos[22480]=1;
cos[22481]=1;
cos[22482]=1;
cos[22483]=1;
cos[22484]=1;
cos[22485]=1;
cos[22486]=1;
cos[22487]=1;
cos[22488]=1;
cos[22489]=1;
cos[22490]=0;
cos[22491]=0;
cos[22492]=0;
cos[22493]=0;
cos[22494]=0;
cos[22495]=0;
cos[22496]=0;
cos[22497]=0;
cos[22498]=0;
cos[22499]=0;
cos[22500]=0;
cos[22501]=0;
cos[22502]=0;
cos[22503]=0;
cos[22504]=0;
cos[22505]=0;
cos[22506]=0;
cos[22507]=0;
cos[22508]=0;
cos[22509]=0;
cos[22510]=0;
cos[22511]=-1;
cos[22512]=-1;
cos[22513]=-1;
cos[22514]=-1;
cos[22515]=-1;
cos[22516]=-1;
cos[22517]=-1;
cos[22518]=-1;
cos[22519]=-1;
cos[22520]=-1;
cos[22521]=-1;
cos[22522]=-1;
cos[22523]=-1;
cos[22524]=-1;
cos[22525]=-1;
cos[22526]=-1;
cos[22527]=-1;
cos[22528]=-1;
cos[22529]=-1;
cos[22530]=-1;
cos[22531]=-2;
cos[22532]=-2;
cos[22533]=-2;
cos[22534]=-2;
cos[22535]=-2;
cos[22536]=-2;
cos[22537]=-2;
cos[22538]=-2;
cos[22539]=-2;
cos[22540]=-2;
cos[22541]=-2;
cos[22542]=-2;
cos[22543]=-2;
cos[22544]=-2;
cos[22545]=-2;
cos[22546]=-2;
cos[22547]=-2;
cos[22548]=-2;
cos[22549]=-2;
cos[22550]=-2;
cos[22551]=-3;
cos[22552]=-3;
cos[22553]=-3;
cos[22554]=-3;
cos[22555]=-3;
cos[22556]=-3;
cos[22557]=-3;
cos[22558]=-3;
cos[22559]=-3;
cos[22560]=-3;
cos[22561]=-3;
cos[22562]=-3;
cos[22563]=-3;
cos[22564]=-3;
cos[22565]=-3;
cos[22566]=-3;
cos[22567]=-3;
cos[22568]=-3;
cos[22569]=-3;
cos[22570]=-3;
cos[22571]=-3;
cos[22572]=-4;
cos[22573]=-4;
cos[22574]=-4;
cos[22575]=-4;
cos[22576]=-4;
cos[22577]=-4;
cos[22578]=-4;
cos[22579]=-4;
cos[22580]=-4;
cos[22581]=-4;
cos[22582]=-4;
cos[22583]=-4;
cos[22584]=-4;
cos[22585]=-4;
cos[22586]=-4;
cos[22587]=-4;
cos[22588]=-4;
cos[22589]=-4;
cos[22590]=-4;
cos[22591]=-4;
cos[22592]=-5;
cos[22593]=-5;
cos[22594]=-5;
cos[22595]=-5;
cos[22596]=-5;
cos[22597]=-5;
cos[22598]=-5;
cos[22599]=-5;
cos[22600]=-5;
cos[22601]=-5;
cos[22602]=-5;
cos[22603]=-5;
cos[22604]=-5;
cos[22605]=-5;
cos[22606]=-5;
cos[22607]=-5;
cos[22608]=-5;
cos[22609]=-5;
cos[22610]=-5;
cos[22611]=-5;
cos[22612]=-5;
cos[22613]=-6;
cos[22614]=-6;
cos[22615]=-6;
cos[22616]=-6;
cos[22617]=-6;
cos[22618]=-6;
cos[22619]=-6;
cos[22620]=-6;
cos[22621]=-6;
cos[22622]=-6;
cos[22623]=-6;
cos[22624]=-6;
cos[22625]=-6;
cos[22626]=-6;
cos[22627]=-6;
cos[22628]=-6;
cos[22629]=-6;
cos[22630]=-6;
cos[22631]=-6;
cos[22632]=-6;
cos[22633]=-7;
cos[22634]=-7;
cos[22635]=-7;
cos[22636]=-7;
cos[22637]=-7;
cos[22638]=-7;
cos[22639]=-7;
cos[22640]=-7;
cos[22641]=-7;
cos[22642]=-7;
cos[22643]=-7;
cos[22644]=-7;
cos[22645]=-7;
cos[22646]=-7;
cos[22647]=-7;
cos[22648]=-7;
cos[22649]=-7;
cos[22650]=-7;
cos[22651]=-7;
cos[22652]=-7;
cos[22653]=-7;
cos[22654]=-8;
cos[22655]=-8;
cos[22656]=-8;
cos[22657]=-8;
cos[22658]=-8;
cos[22659]=-8;
cos[22660]=-8;
cos[22661]=-8;
cos[22662]=-8;
cos[22663]=-8;
cos[22664]=-8;
cos[22665]=-8;
cos[22666]=-8;
cos[22667]=-8;
cos[22668]=-8;
cos[22669]=-8;
cos[22670]=-8;
cos[22671]=-8;
cos[22672]=-8;
cos[22673]=-8;
cos[22674]=-9;
cos[22675]=-9;
cos[22676]=-9;
cos[22677]=-9;
cos[22678]=-9;
cos[22679]=-9;
cos[22680]=-9;
cos[22681]=-9;
cos[22682]=-9;
cos[22683]=-9;
cos[22684]=-9;
cos[22685]=-9;
cos[22686]=-9;
cos[22687]=-9;
cos[22688]=-9;
cos[22689]=-9;
cos[22690]=-9;
cos[22691]=-9;
cos[22692]=-9;
cos[22693]=-9;
cos[22694]=-9;
cos[22695]=-10;
cos[22696]=-10;
cos[22697]=-10;
cos[22698]=-10;
cos[22699]=-10;
cos[22700]=-10;
cos[22701]=-10;
cos[22702]=-10;
cos[22703]=-10;
cos[22704]=-10;
cos[22705]=-10;
cos[22706]=-10;
cos[22707]=-10;
cos[22708]=-10;
cos[22709]=-10;
cos[22710]=-10;
cos[22711]=-10;
cos[22712]=-10;
cos[22713]=-10;
cos[22714]=-10;
cos[22715]=-11;
cos[22716]=-11;
cos[22717]=-11;
cos[22718]=-11;
cos[22719]=-11;
cos[22720]=-11;
cos[22721]=-11;
cos[22722]=-11;
cos[22723]=-11;
cos[22724]=-11;
cos[22725]=-11;
cos[22726]=-11;
cos[22727]=-11;
cos[22728]=-11;
cos[22729]=-11;
cos[22730]=-11;
cos[22731]=-11;
cos[22732]=-11;
cos[22733]=-11;
cos[22734]=-11;
cos[22735]=-11;
cos[22736]=-12;
cos[22737]=-12;
cos[22738]=-12;
cos[22739]=-12;
cos[22740]=-12;
cos[22741]=-12;
cos[22742]=-12;
cos[22743]=-12;
cos[22744]=-12;
cos[22745]=-12;
cos[22746]=-12;
cos[22747]=-12;
cos[22748]=-12;
cos[22749]=-12;
cos[22750]=-12;
cos[22751]=-12;
cos[22752]=-12;
cos[22753]=-12;
cos[22754]=-12;
cos[22755]=-12;
cos[22756]=-13;
cos[22757]=-13;
cos[22758]=-13;
cos[22759]=-13;
cos[22760]=-13;
cos[22761]=-13;
cos[22762]=-13;
cos[22763]=-13;
cos[22764]=-13;
cos[22765]=-13;
cos[22766]=-13;
cos[22767]=-13;
cos[22768]=-13;
cos[22769]=-13;
cos[22770]=-13;
cos[22771]=-13;
cos[22772]=-13;
cos[22773]=-13;
cos[22774]=-13;
cos[22775]=-13;
cos[22776]=-13;
cos[22777]=-14;
cos[22778]=-14;
cos[22779]=-14;
cos[22780]=-14;
cos[22781]=-14;
cos[22782]=-14;
cos[22783]=-14;
cos[22784]=-14;
cos[22785]=-14;
cos[22786]=-14;
cos[22787]=-14;
cos[22788]=-14;
cos[22789]=-14;
cos[22790]=-14;
cos[22791]=-14;
cos[22792]=-14;
cos[22793]=-14;
cos[22794]=-14;
cos[22795]=-14;
cos[22796]=-14;
cos[22797]=-14;
cos[22798]=-15;
cos[22799]=-15;
cos[22800]=-15;
cos[22801]=-15;
cos[22802]=-15;
cos[22803]=-15;
cos[22804]=-15;
cos[22805]=-15;
cos[22806]=-15;
cos[22807]=-15;
cos[22808]=-15;
cos[22809]=-15;
cos[22810]=-15;
cos[22811]=-15;
cos[22812]=-15;
cos[22813]=-15;
cos[22814]=-15;
cos[22815]=-15;
cos[22816]=-15;
cos[22817]=-15;
cos[22818]=-16;
cos[22819]=-16;
cos[22820]=-16;
cos[22821]=-16;
cos[22822]=-16;
cos[22823]=-16;
cos[22824]=-16;
cos[22825]=-16;
cos[22826]=-16;
cos[22827]=-16;
cos[22828]=-16;
cos[22829]=-16;
cos[22830]=-16;
cos[22831]=-16;
cos[22832]=-16;
cos[22833]=-16;
cos[22834]=-16;
cos[22835]=-16;
cos[22836]=-16;
cos[22837]=-16;
cos[22838]=-16;
cos[22839]=-17;
cos[22840]=-17;
cos[22841]=-17;
cos[22842]=-17;
cos[22843]=-17;
cos[22844]=-17;
cos[22845]=-17;
cos[22846]=-17;
cos[22847]=-17;
cos[22848]=-17;
cos[22849]=-17;
cos[22850]=-17;
cos[22851]=-17;
cos[22852]=-17;
cos[22853]=-17;
cos[22854]=-17;
cos[22855]=-17;
cos[22856]=-17;
cos[22857]=-17;
cos[22858]=-17;
cos[22859]=-17;
cos[22860]=-18;
cos[22861]=-18;
cos[22862]=-18;
cos[22863]=-18;
cos[22864]=-18;
cos[22865]=-18;
cos[22866]=-18;
cos[22867]=-18;
cos[22868]=-18;
cos[22869]=-18;
cos[22870]=-18;
cos[22871]=-18;
cos[22872]=-18;
cos[22873]=-18;
cos[22874]=-18;
cos[22875]=-18;
cos[22876]=-18;
cos[22877]=-18;
cos[22878]=-18;
cos[22879]=-18;
cos[22880]=-18;
cos[22881]=-19;
cos[22882]=-19;
cos[22883]=-19;
cos[22884]=-19;
cos[22885]=-19;
cos[22886]=-19;
cos[22887]=-19;
cos[22888]=-19;
cos[22889]=-19;
cos[22890]=-19;
cos[22891]=-19;
cos[22892]=-19;
cos[22893]=-19;
cos[22894]=-19;
cos[22895]=-19;
cos[22896]=-19;
cos[22897]=-19;
cos[22898]=-19;
cos[22899]=-19;
cos[22900]=-19;
cos[22901]=-19;
cos[22902]=-20;
cos[22903]=-20;
cos[22904]=-20;
cos[22905]=-20;
cos[22906]=-20;
cos[22907]=-20;
cos[22908]=-20;
cos[22909]=-20;
cos[22910]=-20;
cos[22911]=-20;
cos[22912]=-20;
cos[22913]=-20;
cos[22914]=-20;
cos[22915]=-20;
cos[22916]=-20;
cos[22917]=-20;
cos[22918]=-20;
cos[22919]=-20;
cos[22920]=-20;
cos[22921]=-20;
cos[22922]=-20;
cos[22923]=-21;
cos[22924]=-21;
cos[22925]=-21;
cos[22926]=-21;
cos[22927]=-21;
cos[22928]=-21;
cos[22929]=-21;
cos[22930]=-21;
cos[22931]=-21;
cos[22932]=-21;
cos[22933]=-21;
cos[22934]=-21;
cos[22935]=-21;
cos[22936]=-21;
cos[22937]=-21;
cos[22938]=-21;
cos[22939]=-21;
cos[22940]=-21;
cos[22941]=-21;
cos[22942]=-21;
cos[22943]=-21;
cos[22944]=-22;
cos[22945]=-22;
cos[22946]=-22;
cos[22947]=-22;
cos[22948]=-22;
cos[22949]=-22;
cos[22950]=-22;
cos[22951]=-22;
cos[22952]=-22;
cos[22953]=-22;
cos[22954]=-22;
cos[22955]=-22;
cos[22956]=-22;
cos[22957]=-22;
cos[22958]=-22;
cos[22959]=-22;
cos[22960]=-22;
cos[22961]=-22;
cos[22962]=-22;
cos[22963]=-22;
cos[22964]=-22;
cos[22965]=-23;
cos[22966]=-23;
cos[22967]=-23;
cos[22968]=-23;
cos[22969]=-23;
cos[22970]=-23;
cos[22971]=-23;
cos[22972]=-23;
cos[22973]=-23;
cos[22974]=-23;
cos[22975]=-23;
cos[22976]=-23;
cos[22977]=-23;
cos[22978]=-23;
cos[22979]=-23;
cos[22980]=-23;
cos[22981]=-23;
cos[22982]=-23;
cos[22983]=-23;
cos[22984]=-23;
cos[22985]=-23;
cos[22986]=-23;
cos[22987]=-24;
cos[22988]=-24;
cos[22989]=-24;
cos[22990]=-24;
cos[22991]=-24;
cos[22992]=-24;
cos[22993]=-24;
cos[22994]=-24;
cos[22995]=-24;
cos[22996]=-24;
cos[22997]=-24;
cos[22998]=-24;
cos[22999]=-24;
cos[23000]=-24;
cos[23001]=-24;
cos[23002]=-24;
cos[23003]=-24;
cos[23004]=-24;
cos[23005]=-24;
cos[23006]=-24;
cos[23007]=-24;
cos[23008]=-25;
cos[23009]=-25;
cos[23010]=-25;
cos[23011]=-25;
cos[23012]=-25;
cos[23013]=-25;
cos[23014]=-25;
cos[23015]=-25;
cos[23016]=-25;
cos[23017]=-25;
cos[23018]=-25;
cos[23019]=-25;
cos[23020]=-25;
cos[23021]=-25;
cos[23022]=-25;
cos[23023]=-25;
cos[23024]=-25;
cos[23025]=-25;
cos[23026]=-25;
cos[23027]=-25;
cos[23028]=-25;
cos[23029]=-25;
cos[23030]=-26;
cos[23031]=-26;
cos[23032]=-26;
cos[23033]=-26;
cos[23034]=-26;
cos[23035]=-26;
cos[23036]=-26;
cos[23037]=-26;
cos[23038]=-26;
cos[23039]=-26;
cos[23040]=-26;
cos[23041]=-26;
cos[23042]=-26;
cos[23043]=-26;
cos[23044]=-26;
cos[23045]=-26;
cos[23046]=-26;
cos[23047]=-26;
cos[23048]=-26;
cos[23049]=-26;
cos[23050]=-26;
cos[23051]=-27;
cos[23052]=-27;
cos[23053]=-27;
cos[23054]=-27;
cos[23055]=-27;
cos[23056]=-27;
cos[23057]=-27;
cos[23058]=-27;
cos[23059]=-27;
cos[23060]=-27;
cos[23061]=-27;
cos[23062]=-27;
cos[23063]=-27;
cos[23064]=-27;
cos[23065]=-27;
cos[23066]=-27;
cos[23067]=-27;
cos[23068]=-27;
cos[23069]=-27;
cos[23070]=-27;
cos[23071]=-27;
cos[23072]=-27;
cos[23073]=-28;
cos[23074]=-28;
cos[23075]=-28;
cos[23076]=-28;
cos[23077]=-28;
cos[23078]=-28;
cos[23079]=-28;
cos[23080]=-28;
cos[23081]=-28;
cos[23082]=-28;
cos[23083]=-28;
cos[23084]=-28;
cos[23085]=-28;
cos[23086]=-28;
cos[23087]=-28;
cos[23088]=-28;
cos[23089]=-28;
cos[23090]=-28;
cos[23091]=-28;
cos[23092]=-28;
cos[23093]=-28;
cos[23094]=-28;
cos[23095]=-29;
cos[23096]=-29;
cos[23097]=-29;
cos[23098]=-29;
cos[23099]=-29;
cos[23100]=-29;
cos[23101]=-29;
cos[23102]=-29;
cos[23103]=-29;
cos[23104]=-29;
cos[23105]=-29;
cos[23106]=-29;
cos[23107]=-29;
cos[23108]=-29;
cos[23109]=-29;
cos[23110]=-29;
cos[23111]=-29;
cos[23112]=-29;
cos[23113]=-29;
cos[23114]=-29;
cos[23115]=-29;
cos[23116]=-29;
cos[23117]=-30;
cos[23118]=-30;
cos[23119]=-30;
cos[23120]=-30;
cos[23121]=-30;
cos[23122]=-30;
cos[23123]=-30;
cos[23124]=-30;
cos[23125]=-30;
cos[23126]=-30;
cos[23127]=-30;
cos[23128]=-30;
cos[23129]=-30;
cos[23130]=-30;
cos[23131]=-30;
cos[23132]=-30;
cos[23133]=-30;
cos[23134]=-30;
cos[23135]=-30;
cos[23136]=-30;
cos[23137]=-30;
cos[23138]=-30;
cos[23139]=-31;
cos[23140]=-31;
cos[23141]=-31;
cos[23142]=-31;
cos[23143]=-31;
cos[23144]=-31;
cos[23145]=-31;
cos[23146]=-31;
cos[23147]=-31;
cos[23148]=-31;
cos[23149]=-31;
cos[23150]=-31;
cos[23151]=-31;
cos[23152]=-31;
cos[23153]=-31;
cos[23154]=-31;
cos[23155]=-31;
cos[23156]=-31;
cos[23157]=-31;
cos[23158]=-31;
cos[23159]=-31;
cos[23160]=-31;
cos[23161]=-32;
cos[23162]=-32;
cos[23163]=-32;
cos[23164]=-32;
cos[23165]=-32;
cos[23166]=-32;
cos[23167]=-32;
cos[23168]=-32;
cos[23169]=-32;
cos[23170]=-32;
cos[23171]=-32;
cos[23172]=-32;
cos[23173]=-32;
cos[23174]=-32;
cos[23175]=-32;
cos[23176]=-32;
cos[23177]=-32;
cos[23178]=-32;
cos[23179]=-32;
cos[23180]=-32;
cos[23181]=-32;
cos[23182]=-32;
cos[23183]=-33;
cos[23184]=-33;
cos[23185]=-33;
cos[23186]=-33;
cos[23187]=-33;
cos[23188]=-33;
cos[23189]=-33;
cos[23190]=-33;
cos[23191]=-33;
cos[23192]=-33;
cos[23193]=-33;
cos[23194]=-33;
cos[23195]=-33;
cos[23196]=-33;
cos[23197]=-33;
cos[23198]=-33;
cos[23199]=-33;
cos[23200]=-33;
cos[23201]=-33;
cos[23202]=-33;
cos[23203]=-33;
cos[23204]=-33;
cos[23205]=-33;
cos[23206]=-34;
cos[23207]=-34;
cos[23208]=-34;
cos[23209]=-34;
cos[23210]=-34;
cos[23211]=-34;
cos[23212]=-34;
cos[23213]=-34;
cos[23214]=-34;
cos[23215]=-34;
cos[23216]=-34;
cos[23217]=-34;
cos[23218]=-34;
cos[23219]=-34;
cos[23220]=-34;
cos[23221]=-34;
cos[23222]=-34;
cos[23223]=-34;
cos[23224]=-34;
cos[23225]=-34;
cos[23226]=-34;
cos[23227]=-34;
cos[23228]=-35;
cos[23229]=-35;
cos[23230]=-35;
cos[23231]=-35;
cos[23232]=-35;
cos[23233]=-35;
cos[23234]=-35;
cos[23235]=-35;
cos[23236]=-35;
cos[23237]=-35;
cos[23238]=-35;
cos[23239]=-35;
cos[23240]=-35;
cos[23241]=-35;
cos[23242]=-35;
cos[23243]=-35;
cos[23244]=-35;
cos[23245]=-35;
cos[23246]=-35;
cos[23247]=-35;
cos[23248]=-35;
cos[23249]=-35;
cos[23250]=-35;
cos[23251]=-36;
cos[23252]=-36;
cos[23253]=-36;
cos[23254]=-36;
cos[23255]=-36;
cos[23256]=-36;
cos[23257]=-36;
cos[23258]=-36;
cos[23259]=-36;
cos[23260]=-36;
cos[23261]=-36;
cos[23262]=-36;
cos[23263]=-36;
cos[23264]=-36;
cos[23265]=-36;
cos[23266]=-36;
cos[23267]=-36;
cos[23268]=-36;
cos[23269]=-36;
cos[23270]=-36;
cos[23271]=-36;
cos[23272]=-36;
cos[23273]=-36;
cos[23274]=-37;
cos[23275]=-37;
cos[23276]=-37;
cos[23277]=-37;
cos[23278]=-37;
cos[23279]=-37;
cos[23280]=-37;
cos[23281]=-37;
cos[23282]=-37;
cos[23283]=-37;
cos[23284]=-37;
cos[23285]=-37;
cos[23286]=-37;
cos[23287]=-37;
cos[23288]=-37;
cos[23289]=-37;
cos[23290]=-37;
cos[23291]=-37;
cos[23292]=-37;
cos[23293]=-37;
cos[23294]=-37;
cos[23295]=-37;
cos[23296]=-37;
cos[23297]=-38;
cos[23298]=-38;
cos[23299]=-38;
cos[23300]=-38;
cos[23301]=-38;
cos[23302]=-38;
cos[23303]=-38;
cos[23304]=-38;
cos[23305]=-38;
cos[23306]=-38;
cos[23307]=-38;
cos[23308]=-38;
cos[23309]=-38;
cos[23310]=-38;
cos[23311]=-38;
cos[23312]=-38;
cos[23313]=-38;
cos[23314]=-38;
cos[23315]=-38;
cos[23316]=-38;
cos[23317]=-38;
cos[23318]=-38;
cos[23319]=-38;
cos[23320]=-38;
cos[23321]=-39;
cos[23322]=-39;
cos[23323]=-39;
cos[23324]=-39;
cos[23325]=-39;
cos[23326]=-39;
cos[23327]=-39;
cos[23328]=-39;
cos[23329]=-39;
cos[23330]=-39;
cos[23331]=-39;
cos[23332]=-39;
cos[23333]=-39;
cos[23334]=-39;
cos[23335]=-39;
cos[23336]=-39;
cos[23337]=-39;
cos[23338]=-39;
cos[23339]=-39;
cos[23340]=-39;
cos[23341]=-39;
cos[23342]=-39;
cos[23343]=-39;
cos[23344]=-40;
cos[23345]=-40;
cos[23346]=-40;
cos[23347]=-40;
cos[23348]=-40;
cos[23349]=-40;
cos[23350]=-40;
cos[23351]=-40;
cos[23352]=-40;
cos[23353]=-40;
cos[23354]=-40;
cos[23355]=-40;
cos[23356]=-40;
cos[23357]=-40;
cos[23358]=-40;
cos[23359]=-40;
cos[23360]=-40;
cos[23361]=-40;
cos[23362]=-40;
cos[23363]=-40;
cos[23364]=-40;
cos[23365]=-40;
cos[23366]=-40;
cos[23367]=-40;
cos[23368]=-41;
cos[23369]=-41;
cos[23370]=-41;
cos[23371]=-41;
cos[23372]=-41;
cos[23373]=-41;
cos[23374]=-41;
cos[23375]=-41;
cos[23376]=-41;
cos[23377]=-41;
cos[23378]=-41;
cos[23379]=-41;
cos[23380]=-41;
cos[23381]=-41;
cos[23382]=-41;
cos[23383]=-41;
cos[23384]=-41;
cos[23385]=-41;
cos[23386]=-41;
cos[23387]=-41;
cos[23388]=-41;
cos[23389]=-41;
cos[23390]=-41;
cos[23391]=-41;
cos[23392]=-42;
cos[23393]=-42;
cos[23394]=-42;
cos[23395]=-42;
cos[23396]=-42;
cos[23397]=-42;
cos[23398]=-42;
cos[23399]=-42;
cos[23400]=-42;
cos[23401]=-42;
cos[23402]=-42;
cos[23403]=-42;
cos[23404]=-42;
cos[23405]=-42;
cos[23406]=-42;
cos[23407]=-42;
cos[23408]=-42;
cos[23409]=-42;
cos[23410]=-42;
cos[23411]=-42;
cos[23412]=-42;
cos[23413]=-42;
cos[23414]=-42;
cos[23415]=-42;
cos[23416]=-43;
cos[23417]=-43;
cos[23418]=-43;
cos[23419]=-43;
cos[23420]=-43;
cos[23421]=-43;
cos[23422]=-43;
cos[23423]=-43;
cos[23424]=-43;
cos[23425]=-43;
cos[23426]=-43;
cos[23427]=-43;
cos[23428]=-43;
cos[23429]=-43;
cos[23430]=-43;
cos[23431]=-43;
cos[23432]=-43;
cos[23433]=-43;
cos[23434]=-43;
cos[23435]=-43;
cos[23436]=-43;
cos[23437]=-43;
cos[23438]=-43;
cos[23439]=-43;
cos[23440]=-44;
cos[23441]=-44;
cos[23442]=-44;
cos[23443]=-44;
cos[23444]=-44;
cos[23445]=-44;
cos[23446]=-44;
cos[23447]=-44;
cos[23448]=-44;
cos[23449]=-44;
cos[23450]=-44;
cos[23451]=-44;
cos[23452]=-44;
cos[23453]=-44;
cos[23454]=-44;
cos[23455]=-44;
cos[23456]=-44;
cos[23457]=-44;
cos[23458]=-44;
cos[23459]=-44;
cos[23460]=-44;
cos[23461]=-44;
cos[23462]=-44;
cos[23463]=-44;
cos[23464]=-44;
cos[23465]=-45;
cos[23466]=-45;
cos[23467]=-45;
cos[23468]=-45;
cos[23469]=-45;
cos[23470]=-45;
cos[23471]=-45;
cos[23472]=-45;
cos[23473]=-45;
cos[23474]=-45;
cos[23475]=-45;
cos[23476]=-45;
cos[23477]=-45;
cos[23478]=-45;
cos[23479]=-45;
cos[23480]=-45;
cos[23481]=-45;
cos[23482]=-45;
cos[23483]=-45;
cos[23484]=-45;
cos[23485]=-45;
cos[23486]=-45;
cos[23487]=-45;
cos[23488]=-45;
cos[23489]=-45;
cos[23490]=-46;
cos[23491]=-46;
cos[23492]=-46;
cos[23493]=-46;
cos[23494]=-46;
cos[23495]=-46;
cos[23496]=-46;
cos[23497]=-46;
cos[23498]=-46;
cos[23499]=-46;
cos[23500]=-46;
cos[23501]=-46;
cos[23502]=-46;
cos[23503]=-46;
cos[23504]=-46;
cos[23505]=-46;
cos[23506]=-46;
cos[23507]=-46;
cos[23508]=-46;
cos[23509]=-46;
cos[23510]=-46;
cos[23511]=-46;
cos[23512]=-46;
cos[23513]=-46;
cos[23514]=-46;
cos[23515]=-47;
cos[23516]=-47;
cos[23517]=-47;
cos[23518]=-47;
cos[23519]=-47;
cos[23520]=-47;
cos[23521]=-47;
cos[23522]=-47;
cos[23523]=-47;
cos[23524]=-47;
cos[23525]=-47;
cos[23526]=-47;
cos[23527]=-47;
cos[23528]=-47;
cos[23529]=-47;
cos[23530]=-47;
cos[23531]=-47;
cos[23532]=-47;
cos[23533]=-47;
cos[23534]=-47;
cos[23535]=-47;
cos[23536]=-47;
cos[23537]=-47;
cos[23538]=-47;
cos[23539]=-47;
cos[23540]=-47;
cos[23541]=-48;
cos[23542]=-48;
cos[23543]=-48;
cos[23544]=-48;
cos[23545]=-48;
cos[23546]=-48;
cos[23547]=-48;
cos[23548]=-48;
cos[23549]=-48;
cos[23550]=-48;
cos[23551]=-48;
cos[23552]=-48;
cos[23553]=-48;
cos[23554]=-48;
cos[23555]=-48;
cos[23556]=-48;
cos[23557]=-48;
cos[23558]=-48;
cos[23559]=-48;
cos[23560]=-48;
cos[23561]=-48;
cos[23562]=-48;
cos[23563]=-48;
cos[23564]=-48;
cos[23565]=-48;
cos[23566]=-49;
cos[23567]=-49;
cos[23568]=-49;
cos[23569]=-49;
cos[23570]=-49;
cos[23571]=-49;
cos[23572]=-49;
cos[23573]=-49;
cos[23574]=-49;
cos[23575]=-49;
cos[23576]=-49;
cos[23577]=-49;
cos[23578]=-49;
cos[23579]=-49;
cos[23580]=-49;
cos[23581]=-49;
cos[23582]=-49;
cos[23583]=-49;
cos[23584]=-49;
cos[23585]=-49;
cos[23586]=-49;
cos[23587]=-49;
cos[23588]=-49;
cos[23589]=-49;
cos[23590]=-49;
cos[23591]=-49;
cos[23592]=-49;
cos[23593]=-50;
cos[23594]=-50;
cos[23595]=-50;
cos[23596]=-50;
cos[23597]=-50;
cos[23598]=-50;
cos[23599]=-50;
cos[23600]=-50;
cos[23601]=-50;
cos[23602]=-50;
cos[23603]=-50;
cos[23604]=-50;
cos[23605]=-50;
cos[23606]=-50;
cos[23607]=-50;
cos[23608]=-50;
cos[23609]=-50;
cos[23610]=-50;
cos[23611]=-50;
cos[23612]=-50;
cos[23613]=-50;
cos[23614]=-50;
cos[23615]=-50;
cos[23616]=-50;
cos[23617]=-50;
cos[23618]=-50;
cos[23619]=-51;
cos[23620]=-51;
cos[23621]=-51;
cos[23622]=-51;
cos[23623]=-51;
cos[23624]=-51;
cos[23625]=-51;
cos[23626]=-51;
cos[23627]=-51;
cos[23628]=-51;
cos[23629]=-51;
cos[23630]=-51;
cos[23631]=-51;
cos[23632]=-51;
cos[23633]=-51;
cos[23634]=-51;
cos[23635]=-51;
cos[23636]=-51;
cos[23637]=-51;
cos[23638]=-51;
cos[23639]=-51;
cos[23640]=-51;
cos[23641]=-51;
cos[23642]=-51;
cos[23643]=-51;
cos[23644]=-51;
cos[23645]=-51;
cos[23646]=-52;
cos[23647]=-52;
cos[23648]=-52;
cos[23649]=-52;
cos[23650]=-52;
cos[23651]=-52;
cos[23652]=-52;
cos[23653]=-52;
cos[23654]=-52;
cos[23655]=-52;
cos[23656]=-52;
cos[23657]=-52;
cos[23658]=-52;
cos[23659]=-52;
cos[23660]=-52;
cos[23661]=-52;
cos[23662]=-52;
cos[23663]=-52;
cos[23664]=-52;
cos[23665]=-52;
cos[23666]=-52;
cos[23667]=-52;
cos[23668]=-52;
cos[23669]=-52;
cos[23670]=-52;
cos[23671]=-52;
cos[23672]=-52;
cos[23673]=-53;
cos[23674]=-53;
cos[23675]=-53;
cos[23676]=-53;
cos[23677]=-53;
cos[23678]=-53;
cos[23679]=-53;
cos[23680]=-53;
cos[23681]=-53;
cos[23682]=-53;
cos[23683]=-53;
cos[23684]=-53;
cos[23685]=-53;
cos[23686]=-53;
cos[23687]=-53;
cos[23688]=-53;
cos[23689]=-53;
cos[23690]=-53;
cos[23691]=-53;
cos[23692]=-53;
cos[23693]=-53;
cos[23694]=-53;
cos[23695]=-53;
cos[23696]=-53;
cos[23697]=-53;
cos[23698]=-53;
cos[23699]=-53;
cos[23700]=-53;
cos[23701]=-54;
cos[23702]=-54;
cos[23703]=-54;
cos[23704]=-54;
cos[23705]=-54;
cos[23706]=-54;
cos[23707]=-54;
cos[23708]=-54;
cos[23709]=-54;
cos[23710]=-54;
cos[23711]=-54;
cos[23712]=-54;
cos[23713]=-54;
cos[23714]=-54;
cos[23715]=-54;
cos[23716]=-54;
cos[23717]=-54;
cos[23718]=-54;
cos[23719]=-54;
cos[23720]=-54;
cos[23721]=-54;
cos[23722]=-54;
cos[23723]=-54;
cos[23724]=-54;
cos[23725]=-54;
cos[23726]=-54;
cos[23727]=-54;
cos[23728]=-54;
cos[23729]=-55;
cos[23730]=-55;
cos[23731]=-55;
cos[23732]=-55;
cos[23733]=-55;
cos[23734]=-55;
cos[23735]=-55;
cos[23736]=-55;
cos[23737]=-55;
cos[23738]=-55;
cos[23739]=-55;
cos[23740]=-55;
cos[23741]=-55;
cos[23742]=-55;
cos[23743]=-55;
cos[23744]=-55;
cos[23745]=-55;
cos[23746]=-55;
cos[23747]=-55;
cos[23748]=-55;
cos[23749]=-55;
cos[23750]=-55;
cos[23751]=-55;
cos[23752]=-55;
cos[23753]=-55;
cos[23754]=-55;
cos[23755]=-55;
cos[23756]=-55;
cos[23757]=-55;
cos[23758]=-56;
cos[23759]=-56;
cos[23760]=-56;
cos[23761]=-56;
cos[23762]=-56;
cos[23763]=-56;
cos[23764]=-56;
cos[23765]=-56;
cos[23766]=-56;
cos[23767]=-56;
cos[23768]=-56;
cos[23769]=-56;
cos[23770]=-56;
cos[23771]=-56;
cos[23772]=-56;
cos[23773]=-56;
cos[23774]=-56;
cos[23775]=-56;
cos[23776]=-56;
cos[23777]=-56;
cos[23778]=-56;
cos[23779]=-56;
cos[23780]=-56;
cos[23781]=-56;
cos[23782]=-56;
cos[23783]=-56;
cos[23784]=-56;
cos[23785]=-56;
cos[23786]=-56;
cos[23787]=-57;
cos[23788]=-57;
cos[23789]=-57;
cos[23790]=-57;
cos[23791]=-57;
cos[23792]=-57;
cos[23793]=-57;
cos[23794]=-57;
cos[23795]=-57;
cos[23796]=-57;
cos[23797]=-57;
cos[23798]=-57;
cos[23799]=-57;
cos[23800]=-57;
cos[23801]=-57;
cos[23802]=-57;
cos[23803]=-57;
cos[23804]=-57;
cos[23805]=-57;
cos[23806]=-57;
cos[23807]=-57;
cos[23808]=-57;
cos[23809]=-57;
cos[23810]=-57;
cos[23811]=-57;
cos[23812]=-57;
cos[23813]=-57;
cos[23814]=-57;
cos[23815]=-57;
cos[23816]=-57;
cos[23817]=-58;
cos[23818]=-58;
cos[23819]=-58;
cos[23820]=-58;
cos[23821]=-58;
cos[23822]=-58;
cos[23823]=-58;
cos[23824]=-58;
cos[23825]=-58;
cos[23826]=-58;
cos[23827]=-58;
cos[23828]=-58;
cos[23829]=-58;
cos[23830]=-58;
cos[23831]=-58;
cos[23832]=-58;
cos[23833]=-58;
cos[23834]=-58;
cos[23835]=-58;
cos[23836]=-58;
cos[23837]=-58;
cos[23838]=-58;
cos[23839]=-58;
cos[23840]=-58;
cos[23841]=-58;
cos[23842]=-58;
cos[23843]=-58;
cos[23844]=-58;
cos[23845]=-58;
cos[23846]=-58;
cos[23847]=-59;
cos[23848]=-59;
cos[23849]=-59;
cos[23850]=-59;
cos[23851]=-59;
cos[23852]=-59;
cos[23853]=-59;
cos[23854]=-59;
cos[23855]=-59;
cos[23856]=-59;
cos[23857]=-59;
cos[23858]=-59;
cos[23859]=-59;
cos[23860]=-59;
cos[23861]=-59;
cos[23862]=-59;
cos[23863]=-59;
cos[23864]=-59;
cos[23865]=-59;
cos[23866]=-59;
cos[23867]=-59;
cos[23868]=-59;
cos[23869]=-59;
cos[23870]=-59;
cos[23871]=-59;
cos[23872]=-59;
cos[23873]=-59;
cos[23874]=-59;
cos[23875]=-59;
cos[23876]=-59;
cos[23877]=-59;
cos[23878]=-60;
cos[23879]=-60;
cos[23880]=-60;
cos[23881]=-60;
cos[23882]=-60;
cos[23883]=-60;
cos[23884]=-60;
cos[23885]=-60;
cos[23886]=-60;
cos[23887]=-60;
cos[23888]=-60;
cos[23889]=-60;
cos[23890]=-60;
cos[23891]=-60;
cos[23892]=-60;
cos[23893]=-60;
cos[23894]=-60;
cos[23895]=-60;
cos[23896]=-60;
cos[23897]=-60;
cos[23898]=-60;
cos[23899]=-60;
cos[23900]=-60;
cos[23901]=-60;
cos[23902]=-60;
cos[23903]=-60;
cos[23904]=-60;
cos[23905]=-60;
cos[23906]=-60;
cos[23907]=-60;
cos[23908]=-60;
cos[23909]=-60;
cos[23910]=-61;
cos[23911]=-61;
cos[23912]=-61;
cos[23913]=-61;
cos[23914]=-61;
cos[23915]=-61;
cos[23916]=-61;
cos[23917]=-61;
cos[23918]=-61;
cos[23919]=-61;
cos[23920]=-61;
cos[23921]=-61;
cos[23922]=-61;
cos[23923]=-61;
cos[23924]=-61;
cos[23925]=-61;
cos[23926]=-61;
cos[23927]=-61;
cos[23928]=-61;
cos[23929]=-61;
cos[23930]=-61;
cos[23931]=-61;
cos[23932]=-61;
cos[23933]=-61;
cos[23934]=-61;
cos[23935]=-61;
cos[23936]=-61;
cos[23937]=-61;
cos[23938]=-61;
cos[23939]=-61;
cos[23940]=-61;
cos[23941]=-61;
cos[23942]=-61;
cos[23943]=-62;
cos[23944]=-62;
cos[23945]=-62;
cos[23946]=-62;
cos[23947]=-62;
cos[23948]=-62;
cos[23949]=-62;
cos[23950]=-62;
cos[23951]=-62;
cos[23952]=-62;
cos[23953]=-62;
cos[23954]=-62;
cos[23955]=-62;
cos[23956]=-62;
cos[23957]=-62;
cos[23958]=-62;
cos[23959]=-62;
cos[23960]=-62;
cos[23961]=-62;
cos[23962]=-62;
cos[23963]=-62;
cos[23964]=-62;
cos[23965]=-62;
cos[23966]=-62;
cos[23967]=-62;
cos[23968]=-62;
cos[23969]=-62;
cos[23970]=-62;
cos[23971]=-62;
cos[23972]=-62;
cos[23973]=-62;
cos[23974]=-62;
cos[23975]=-62;
cos[23976]=-63;
cos[23977]=-63;
cos[23978]=-63;
cos[23979]=-63;
cos[23980]=-63;
cos[23981]=-63;
cos[23982]=-63;
cos[23983]=-63;
cos[23984]=-63;
cos[23985]=-63;
cos[23986]=-63;
cos[23987]=-63;
cos[23988]=-63;
cos[23989]=-63;
cos[23990]=-63;
cos[23991]=-63;
cos[23992]=-63;
cos[23993]=-63;
cos[23994]=-63;
cos[23995]=-63;
cos[23996]=-63;
cos[23997]=-63;
cos[23998]=-63;
cos[23999]=-63;
cos[24000]=-63;
cos[24001]=-63;
cos[24002]=-63;
cos[24003]=-63;
cos[24004]=-63;
cos[24005]=-63;
cos[24006]=-63;
cos[24007]=-63;
cos[24008]=-63;
cos[24009]=-63;
cos[24010]=-63;
cos[24011]=-64;
cos[24012]=-64;
cos[24013]=-64;
cos[24014]=-64;
cos[24015]=-64;
cos[24016]=-64;
cos[24017]=-64;
cos[24018]=-64;
cos[24019]=-64;
cos[24020]=-64;
cos[24021]=-64;
cos[24022]=-64;
cos[24023]=-64;
cos[24024]=-64;
cos[24025]=-64;
cos[24026]=-64;
cos[24027]=-64;
cos[24028]=-64;
cos[24029]=-64;
cos[24030]=-64;
cos[24031]=-64;
cos[24032]=-64;
cos[24033]=-64;
cos[24034]=-64;
cos[24035]=-64;
cos[24036]=-64;
cos[24037]=-64;
cos[24038]=-64;
cos[24039]=-64;
cos[24040]=-64;
cos[24041]=-64;
cos[24042]=-64;
cos[24043]=-64;
cos[24044]=-64;
cos[24045]=-64;
cos[24046]=-65;
cos[24047]=-65;
cos[24048]=-65;
cos[24049]=-65;
cos[24050]=-65;
cos[24051]=-65;
cos[24052]=-65;
cos[24053]=-65;
cos[24054]=-65;
cos[24055]=-65;
cos[24056]=-65;
cos[24057]=-65;
cos[24058]=-65;
cos[24059]=-65;
cos[24060]=-65;
cos[24061]=-65;
cos[24062]=-65;
cos[24063]=-65;
cos[24064]=-65;
cos[24065]=-65;
cos[24066]=-65;
cos[24067]=-65;
cos[24068]=-65;
cos[24069]=-65;
cos[24070]=-65;
cos[24071]=-65;
cos[24072]=-65;
cos[24073]=-65;
cos[24074]=-65;
cos[24075]=-65;
cos[24076]=-65;
cos[24077]=-65;
cos[24078]=-65;
cos[24079]=-65;
cos[24080]=-65;
cos[24081]=-65;
cos[24082]=-65;
cos[24083]=-66;
cos[24084]=-66;
cos[24085]=-66;
cos[24086]=-66;
cos[24087]=-66;
cos[24088]=-66;
cos[24089]=-66;
cos[24090]=-66;
cos[24091]=-66;
cos[24092]=-66;
cos[24093]=-66;
cos[24094]=-66;
cos[24095]=-66;
cos[24096]=-66;
cos[24097]=-66;
cos[24098]=-66;
cos[24099]=-66;
cos[24100]=-66;
cos[24101]=-66;
cos[24102]=-66;
cos[24103]=-66;
cos[24104]=-66;
cos[24105]=-66;
cos[24106]=-66;
cos[24107]=-66;
cos[24108]=-66;
cos[24109]=-66;
cos[24110]=-66;
cos[24111]=-66;
cos[24112]=-66;
cos[24113]=-66;
cos[24114]=-66;
cos[24115]=-66;
cos[24116]=-66;
cos[24117]=-66;
cos[24118]=-66;
cos[24119]=-66;
cos[24120]=-66;
cos[24121]=-67;
cos[24122]=-67;
cos[24123]=-67;
cos[24124]=-67;
cos[24125]=-67;
cos[24126]=-67;
cos[24127]=-67;
cos[24128]=-67;
cos[24129]=-67;
cos[24130]=-67;
cos[24131]=-67;
cos[24132]=-67;
cos[24133]=-67;
cos[24134]=-67;
cos[24135]=-67;
cos[24136]=-67;
cos[24137]=-67;
cos[24138]=-67;
cos[24139]=-67;
cos[24140]=-67;
cos[24141]=-67;
cos[24142]=-67;
cos[24143]=-67;
cos[24144]=-67;
cos[24145]=-67;
cos[24146]=-67;
cos[24147]=-67;
cos[24148]=-67;
cos[24149]=-67;
cos[24150]=-67;
cos[24151]=-67;
cos[24152]=-67;
cos[24153]=-67;
cos[24154]=-67;
cos[24155]=-67;
cos[24156]=-67;
cos[24157]=-67;
cos[24158]=-67;
cos[24159]=-67;
cos[24160]=-67;
cos[24161]=-68;
cos[24162]=-68;
cos[24163]=-68;
cos[24164]=-68;
cos[24165]=-68;
cos[24166]=-68;
cos[24167]=-68;
cos[24168]=-68;
cos[24169]=-68;
cos[24170]=-68;
cos[24171]=-68;
cos[24172]=-68;
cos[24173]=-68;
cos[24174]=-68;
cos[24175]=-68;
cos[24176]=-68;
cos[24177]=-68;
cos[24178]=-68;
cos[24179]=-68;
cos[24180]=-68;
cos[24181]=-68;
cos[24182]=-68;
cos[24183]=-68;
cos[24184]=-68;
cos[24185]=-68;
cos[24186]=-68;
cos[24187]=-68;
cos[24188]=-68;
cos[24189]=-68;
cos[24190]=-68;
cos[24191]=-68;
cos[24192]=-68;
cos[24193]=-68;
cos[24194]=-68;
cos[24195]=-68;
cos[24196]=-68;
cos[24197]=-68;
cos[24198]=-68;
cos[24199]=-68;
cos[24200]=-68;
cos[24201]=-68;
cos[24202]=-69;
cos[24203]=-69;
cos[24204]=-69;
cos[24205]=-69;
cos[24206]=-69;
cos[24207]=-69;
cos[24208]=-69;
cos[24209]=-69;
cos[24210]=-69;
cos[24211]=-69;
cos[24212]=-69;
cos[24213]=-69;
cos[24214]=-69;
cos[24215]=-69;
cos[24216]=-69;
cos[24217]=-69;
cos[24218]=-69;
cos[24219]=-69;
cos[24220]=-69;
cos[24221]=-69;
cos[24222]=-69;
cos[24223]=-69;
cos[24224]=-69;
cos[24225]=-69;
cos[24226]=-69;
cos[24227]=-69;
cos[24228]=-69;
cos[24229]=-69;
cos[24230]=-69;
cos[24231]=-69;
cos[24232]=-69;
cos[24233]=-69;
cos[24234]=-69;
cos[24235]=-69;
cos[24236]=-69;
cos[24237]=-69;
cos[24238]=-69;
cos[24239]=-69;
cos[24240]=-69;
cos[24241]=-69;
cos[24242]=-69;
cos[24243]=-69;
cos[24244]=-69;
cos[24245]=-69;
cos[24246]=-70;
cos[24247]=-70;
cos[24248]=-70;
cos[24249]=-70;
cos[24250]=-70;
cos[24251]=-70;
cos[24252]=-70;
cos[24253]=-70;
cos[24254]=-70;
cos[24255]=-70;
cos[24256]=-70;
cos[24257]=-70;
cos[24258]=-70;
cos[24259]=-70;
cos[24260]=-70;
cos[24261]=-70;
cos[24262]=-70;
cos[24263]=-70;
cos[24264]=-70;
cos[24265]=-70;
cos[24266]=-70;
cos[24267]=-70;
cos[24268]=-70;
cos[24269]=-70;
cos[24270]=-70;
cos[24271]=-70;
cos[24272]=-70;
cos[24273]=-70;
cos[24274]=-70;
cos[24275]=-70;
cos[24276]=-70;
cos[24277]=-70;
cos[24278]=-70;
cos[24279]=-70;
cos[24280]=-70;
cos[24281]=-70;
cos[24282]=-70;
cos[24283]=-70;
cos[24284]=-70;
cos[24285]=-70;
cos[24286]=-70;
cos[24287]=-70;
cos[24288]=-70;
cos[24289]=-70;
cos[24290]=-70;
cos[24291]=-71;
cos[24292]=-71;
cos[24293]=-71;
cos[24294]=-71;
cos[24295]=-71;
cos[24296]=-71;
cos[24297]=-71;
cos[24298]=-71;
cos[24299]=-71;
cos[24300]=-71;
cos[24301]=-71;
cos[24302]=-71;
cos[24303]=-71;
cos[24304]=-71;
cos[24305]=-71;
cos[24306]=-71;
cos[24307]=-71;
cos[24308]=-71;
cos[24309]=-71;
cos[24310]=-71;
cos[24311]=-71;
cos[24312]=-71;
cos[24313]=-71;
cos[24314]=-71;
cos[24315]=-71;
cos[24316]=-71;
cos[24317]=-71;
cos[24318]=-71;
cos[24319]=-71;
cos[24320]=-71;
cos[24321]=-71;
cos[24322]=-71;
cos[24323]=-71;
cos[24324]=-71;
cos[24325]=-71;
cos[24326]=-71;
cos[24327]=-71;
cos[24328]=-71;
cos[24329]=-71;
cos[24330]=-71;
cos[24331]=-71;
cos[24332]=-71;
cos[24333]=-71;
cos[24334]=-71;
cos[24335]=-71;
cos[24336]=-71;
cos[24337]=-71;
cos[24338]=-71;
cos[24339]=-71;
cos[24340]=-72;
cos[24341]=-72;
cos[24342]=-72;
cos[24343]=-72;
cos[24344]=-72;
cos[24345]=-72;
cos[24346]=-72;
cos[24347]=-72;
cos[24348]=-72;
cos[24349]=-72;
cos[24350]=-72;
cos[24351]=-72;
cos[24352]=-72;
cos[24353]=-72;
cos[24354]=-72;
cos[24355]=-72;
cos[24356]=-72;
cos[24357]=-72;
cos[24358]=-72;
cos[24359]=-72;
cos[24360]=-72;
cos[24361]=-72;
cos[24362]=-72;
cos[24363]=-72;
cos[24364]=-72;
cos[24365]=-72;
cos[24366]=-72;
cos[24367]=-72;
cos[24368]=-72;
cos[24369]=-72;
cos[24370]=-72;
cos[24371]=-72;
cos[24372]=-72;
cos[24373]=-72;
cos[24374]=-72;
cos[24375]=-72;
cos[24376]=-72;
cos[24377]=-72;
cos[24378]=-72;
cos[24379]=-72;
cos[24380]=-72;
cos[24381]=-72;
cos[24382]=-72;
cos[24383]=-72;
cos[24384]=-72;
cos[24385]=-72;
cos[24386]=-72;
cos[24387]=-72;
cos[24388]=-72;
cos[24389]=-72;
cos[24390]=-72;
cos[24391]=-72;
cos[24392]=-72;
cos[24393]=-73;
cos[24394]=-73;
cos[24395]=-73;
cos[24396]=-73;
cos[24397]=-73;
cos[24398]=-73;
cos[24399]=-73;
cos[24400]=-73;
cos[24401]=-73;
cos[24402]=-73;
cos[24403]=-73;
cos[24404]=-73;
cos[24405]=-73;
cos[24406]=-73;
cos[24407]=-73;
cos[24408]=-73;
cos[24409]=-73;
cos[24410]=-73;
cos[24411]=-73;
cos[24412]=-73;
cos[24413]=-73;
cos[24414]=-73;
cos[24415]=-73;
cos[24416]=-73;
cos[24417]=-73;
cos[24418]=-73;
cos[24419]=-73;
cos[24420]=-73;
cos[24421]=-73;
cos[24422]=-73;
cos[24423]=-73;
cos[24424]=-73;
cos[24425]=-73;
cos[24426]=-73;
cos[24427]=-73;
cos[24428]=-73;
cos[24429]=-73;
cos[24430]=-73;
cos[24431]=-73;
cos[24432]=-73;
cos[24433]=-73;
cos[24434]=-73;
cos[24435]=-73;
cos[24436]=-73;
cos[24437]=-73;
cos[24438]=-73;
cos[24439]=-73;
cos[24440]=-73;
cos[24441]=-73;
cos[24442]=-73;
cos[24443]=-73;
cos[24444]=-73;
cos[24445]=-73;
cos[24446]=-73;
cos[24447]=-73;
cos[24448]=-73;
cos[24449]=-73;
cos[24450]=-74;
cos[24451]=-74;
cos[24452]=-74;
cos[24453]=-74;
cos[24454]=-74;
cos[24455]=-74;
cos[24456]=-74;
cos[24457]=-74;
cos[24458]=-74;
cos[24459]=-74;
cos[24460]=-74;
cos[24461]=-74;
cos[24462]=-74;
cos[24463]=-74;
cos[24464]=-74;
cos[24465]=-74;
cos[24466]=-74;
cos[24467]=-74;
cos[24468]=-74;
cos[24469]=-74;
cos[24470]=-74;
cos[24471]=-74;
cos[24472]=-74;
cos[24473]=-74;
cos[24474]=-74;
cos[24475]=-74;
cos[24476]=-74;
cos[24477]=-74;
cos[24478]=-74;
cos[24479]=-74;
cos[24480]=-74;
cos[24481]=-74;
cos[24482]=-74;
cos[24483]=-74;
cos[24484]=-74;
cos[24485]=-74;
cos[24486]=-74;
cos[24487]=-74;
cos[24488]=-74;
cos[24489]=-74;
cos[24490]=-74;
cos[24491]=-74;
cos[24492]=-74;
cos[24493]=-74;
cos[24494]=-74;
cos[24495]=-74;
cos[24496]=-74;
cos[24497]=-74;
cos[24498]=-74;
cos[24499]=-74;
cos[24500]=-74;
cos[24501]=-74;
cos[24502]=-74;
cos[24503]=-74;
cos[24504]=-74;
cos[24505]=-74;
cos[24506]=-74;
cos[24507]=-74;
cos[24508]=-74;
cos[24509]=-74;
cos[24510]=-74;
cos[24511]=-74;
cos[24512]=-74;
cos[24513]=-74;
cos[24514]=-75;
cos[24515]=-75;
cos[24516]=-75;
cos[24517]=-75;
cos[24518]=-75;
cos[24519]=-75;
cos[24520]=-75;
cos[24521]=-75;
cos[24522]=-75;
cos[24523]=-75;
cos[24524]=-75;
cos[24525]=-75;
cos[24526]=-75;
cos[24527]=-75;
cos[24528]=-75;
cos[24529]=-75;
cos[24530]=-75;
cos[24531]=-75;
cos[24532]=-75;
cos[24533]=-75;
cos[24534]=-75;
cos[24535]=-75;
cos[24536]=-75;
cos[24537]=-75;
cos[24538]=-75;
cos[24539]=-75;
cos[24540]=-75;
cos[24541]=-75;
cos[24542]=-75;
cos[24543]=-75;
cos[24544]=-75;
cos[24545]=-75;
cos[24546]=-75;
cos[24547]=-75;
cos[24548]=-75;
cos[24549]=-75;
cos[24550]=-75;
cos[24551]=-75;
cos[24552]=-75;
cos[24553]=-75;
cos[24554]=-75;
cos[24555]=-75;
cos[24556]=-75;
cos[24557]=-75;
cos[24558]=-75;
cos[24559]=-75;
cos[24560]=-75;
cos[24561]=-75;
cos[24562]=-75;
cos[24563]=-75;
cos[24564]=-75;
cos[24565]=-75;
cos[24566]=-75;
cos[24567]=-75;
cos[24568]=-75;
cos[24569]=-75;
cos[24570]=-75;
cos[24571]=-75;
cos[24572]=-75;
cos[24573]=-75;
cos[24574]=-75;
cos[24575]=-75;
cos[24576]=-75;
cos[24577]=-75;
cos[24578]=-75;
cos[24579]=-75;
cos[24580]=-75;
cos[24581]=-75;
cos[24582]=-75;
cos[24583]=-75;
cos[24584]=-75;
cos[24585]=-75;
cos[24586]=-75;
cos[24587]=-76;
cos[24588]=-76;
cos[24589]=-76;
cos[24590]=-76;
cos[24591]=-76;
cos[24592]=-76;
cos[24593]=-76;
cos[24594]=-76;
cos[24595]=-76;
cos[24596]=-76;
cos[24597]=-76;
cos[24598]=-76;
cos[24599]=-76;
cos[24600]=-76;
cos[24601]=-76;
cos[24602]=-76;
cos[24603]=-76;
cos[24604]=-76;
cos[24605]=-76;
cos[24606]=-76;
cos[24607]=-76;
cos[24608]=-76;
cos[24609]=-76;
cos[24610]=-76;
cos[24611]=-76;
cos[24612]=-76;
cos[24613]=-76;
cos[24614]=-76;
cos[24615]=-76;
cos[24616]=-76;
cos[24617]=-76;
cos[24618]=-76;
cos[24619]=-76;
cos[24620]=-76;
cos[24621]=-76;
cos[24622]=-76;
cos[24623]=-76;
cos[24624]=-76;
cos[24625]=-76;
cos[24626]=-76;
cos[24627]=-76;
cos[24628]=-76;
cos[24629]=-76;
cos[24630]=-76;
cos[24631]=-76;
cos[24632]=-76;
cos[24633]=-76;
cos[24634]=-76;
cos[24635]=-76;
cos[24636]=-76;
cos[24637]=-76;
cos[24638]=-76;
cos[24639]=-76;
cos[24640]=-76;
cos[24641]=-76;
cos[24642]=-76;
cos[24643]=-76;
cos[24644]=-76;
cos[24645]=-76;
cos[24646]=-76;
cos[24647]=-76;
cos[24648]=-76;
cos[24649]=-76;
cos[24650]=-76;
cos[24651]=-76;
cos[24652]=-76;
cos[24653]=-76;
cos[24654]=-76;
cos[24655]=-76;
cos[24656]=-76;
cos[24657]=-76;
cos[24658]=-76;
cos[24659]=-76;
cos[24660]=-76;
cos[24661]=-76;
cos[24662]=-76;
cos[24663]=-76;
cos[24664]=-76;
cos[24665]=-76;
cos[24666]=-76;
cos[24667]=-76;
cos[24668]=-76;
cos[24669]=-76;
cos[24670]=-76;
cos[24671]=-76;
cos[24672]=-76;
cos[24673]=-76;
cos[24674]=-76;
cos[24675]=-77;
cos[24676]=-77;
cos[24677]=-77;
cos[24678]=-77;
cos[24679]=-77;
cos[24680]=-77;
cos[24681]=-77;
cos[24682]=-77;
cos[24683]=-77;
cos[24684]=-77;
cos[24685]=-77;
cos[24686]=-77;
cos[24687]=-77;
cos[24688]=-77;
cos[24689]=-77;
cos[24690]=-77;
cos[24691]=-77;
cos[24692]=-77;
cos[24693]=-77;
cos[24694]=-77;
cos[24695]=-77;
cos[24696]=-77;
cos[24697]=-77;
cos[24698]=-77;
cos[24699]=-77;
cos[24700]=-77;
cos[24701]=-77;
cos[24702]=-77;
cos[24703]=-77;
cos[24704]=-77;
cos[24705]=-77;
cos[24706]=-77;
cos[24707]=-77;
cos[24708]=-77;
cos[24709]=-77;
cos[24710]=-77;
cos[24711]=-77;
cos[24712]=-77;
cos[24713]=-77;
cos[24714]=-77;
cos[24715]=-77;
cos[24716]=-77;
cos[24717]=-77;
cos[24718]=-77;
cos[24719]=-77;
cos[24720]=-77;
cos[24721]=-77;
cos[24722]=-77;
cos[24723]=-77;
cos[24724]=-77;
cos[24725]=-77;
cos[24726]=-77;
cos[24727]=-77;
cos[24728]=-77;
cos[24729]=-77;
cos[24730]=-77;
cos[24731]=-77;
cos[24732]=-77;
cos[24733]=-77;
cos[24734]=-77;
cos[24735]=-77;
cos[24736]=-77;
cos[24737]=-77;
cos[24738]=-77;
cos[24739]=-77;
cos[24740]=-77;
cos[24741]=-77;
cos[24742]=-77;
cos[24743]=-77;
cos[24744]=-77;
cos[24745]=-77;
cos[24746]=-77;
cos[24747]=-77;
cos[24748]=-77;
cos[24749]=-77;
cos[24750]=-77;
cos[24751]=-77;
cos[24752]=-77;
cos[24753]=-77;
cos[24754]=-77;
cos[24755]=-77;
cos[24756]=-77;
cos[24757]=-77;
cos[24758]=-77;
cos[24759]=-77;
cos[24760]=-77;
cos[24761]=-77;
cos[24762]=-77;
cos[24763]=-77;
cos[24764]=-77;
cos[24765]=-77;
cos[24766]=-77;
cos[24767]=-77;
cos[24768]=-77;
cos[24769]=-77;
cos[24770]=-77;
cos[24771]=-77;
cos[24772]=-77;
cos[24773]=-77;
cos[24774]=-77;
cos[24775]=-77;
cos[24776]=-77;
cos[24777]=-77;
cos[24778]=-77;
cos[24779]=-77;
cos[24780]=-77;
cos[24781]=-77;
cos[24782]=-77;
cos[24783]=-77;
cos[24784]=-77;
cos[24785]=-77;
cos[24786]=-77;
cos[24787]=-77;
cos[24788]=-77;
cos[24789]=-77;
cos[24790]=-77;
cos[24791]=-77;
cos[24792]=-77;
cos[24793]=-77;
cos[24794]=-77;
cos[24795]=-77;
cos[24796]=-77;
cos[24797]=-77;
cos[24798]=-77;
cos[24799]=-78;
cos[24800]=-78;
cos[24801]=-78;
cos[24802]=-78;
cos[24803]=-78;
cos[24804]=-78;
cos[24805]=-78;
cos[24806]=-78;
cos[24807]=-78;
cos[24808]=-78;
cos[24809]=-78;
cos[24810]=-78;
cos[24811]=-78;
cos[24812]=-78;
cos[24813]=-78;
cos[24814]=-78;
cos[24815]=-78;
cos[24816]=-78;
cos[24817]=-78;
cos[24818]=-78;
cos[24819]=-78;
cos[24820]=-78;
cos[24821]=-78;
cos[24822]=-78;
cos[24823]=-78;
cos[24824]=-78;
cos[24825]=-78;
cos[24826]=-78;
cos[24827]=-78;
cos[24828]=-78;
cos[24829]=-78;
cos[24830]=-78;
cos[24831]=-78;
cos[24832]=-78;
cos[24833]=-78;
cos[24834]=-78;
cos[24835]=-78;
cos[24836]=-78;
cos[24837]=-78;
cos[24838]=-78;
cos[24839]=-78;
cos[24840]=-78;
cos[24841]=-78;
cos[24842]=-78;
cos[24843]=-78;
cos[24844]=-78;
cos[24845]=-78;
cos[24846]=-78;
cos[24847]=-78;
cos[24848]=-78;
cos[24849]=-78;
cos[24850]=-78;
cos[24851]=-78;
cos[24852]=-78;
cos[24853]=-78;
cos[24854]=-78;
cos[24855]=-78;
cos[24856]=-78;
cos[24857]=-78;
cos[24858]=-78;
cos[24859]=-78;
cos[24860]=-78;
cos[24861]=-78;
cos[24862]=-78;
cos[24863]=-78;
cos[24864]=-78;
cos[24865]=-78;
cos[24866]=-78;
cos[24867]=-78;
cos[24868]=-78;
cos[24869]=-78;
cos[24870]=-78;
cos[24871]=-78;
cos[24872]=-78;
cos[24873]=-78;
cos[24874]=-78;
cos[24875]=-78;
cos[24876]=-78;
cos[24877]=-78;
cos[24878]=-78;
cos[24879]=-78;
cos[24880]=-78;
cos[24881]=-78;
cos[24882]=-78;
cos[24883]=-78;
cos[24884]=-78;
cos[24885]=-78;
cos[24886]=-78;
cos[24887]=-78;
cos[24888]=-78;
cos[24889]=-78;
cos[24890]=-78;
cos[24891]=-78;
cos[24892]=-78;
cos[24893]=-78;
cos[24894]=-78;
cos[24895]=-78;
cos[24896]=-78;
cos[24897]=-78;
cos[24898]=-78;
cos[24899]=-78;
cos[24900]=-78;
cos[24901]=-78;
cos[24902]=-78;
cos[24903]=-78;
cos[24904]=-78;
cos[24905]=-78;
cos[24906]=-78;
cos[24907]=-78;
cos[24908]=-78;
cos[24909]=-78;
cos[24910]=-78;
cos[24911]=-78;
cos[24912]=-78;
cos[24913]=-78;
cos[24914]=-78;
cos[24915]=-78;
cos[24916]=-78;
cos[24917]=-78;
cos[24918]=-78;
cos[24919]=-78;
cos[24920]=-78;
cos[24921]=-78;
cos[24922]=-78;
cos[24923]=-78;
cos[24924]=-78;
cos[24925]=-78;
cos[24926]=-78;
cos[24927]=-78;
cos[24928]=-78;
cos[24929]=-78;
cos[24930]=-78;
cos[24931]=-78;
cos[24932]=-78;
cos[24933]=-78;
cos[24934]=-78;
cos[24935]=-78;
cos[24936]=-78;
cos[24937]=-78;
cos[24938]=-78;
cos[24939]=-78;
cos[24940]=-78;
cos[24941]=-78;
cos[24942]=-78;
cos[24943]=-78;
cos[24944]=-78;
cos[24945]=-78;
cos[24946]=-78;
cos[24947]=-78;
cos[24948]=-78;
cos[24949]=-78;
cos[24950]=-78;
cos[24951]=-78;
cos[24952]=-78;
cos[24953]=-78;
cos[24954]=-78;
cos[24955]=-78;
cos[24956]=-78;
cos[24957]=-78;
cos[24958]=-78;
cos[24959]=-78;
cos[24960]=-78;
cos[24961]=-78;
cos[24962]=-78;
cos[24963]=-78;
cos[24964]=-78;
cos[24965]=-78;
cos[24966]=-78;
cos[24967]=-78;
cos[24968]=-78;
cos[24969]=-78;
cos[24970]=-78;
cos[24971]=-78;
cos[24972]=-78;
cos[24973]=-78;
cos[24974]=-78;
cos[24975]=-78;
cos[24976]=-78;
cos[24977]=-78;
cos[24978]=-78;
cos[24979]=-78;
cos[24980]=-78;
cos[24981]=-78;
cos[24982]=-78;
cos[24983]=-78;
cos[24984]=-78;
cos[24985]=-78;
cos[24986]=-78;
cos[24987]=-78;
cos[24988]=-78;
cos[24989]=-78;
cos[24990]=-78;
cos[24991]=-78;
cos[24992]=-78;
cos[24993]=-78;
cos[24994]=-78;
cos[24995]=-78;
cos[24996]=-78;
cos[24997]=-78;
cos[24998]=-78;
cos[24999]=-78;
cos[25000]=-78;
cos[25001]=-78;
cos[25002]=-78;
cos[25003]=-78;
cos[25004]=-78;
cos[25005]=-78;
cos[25006]=-78;
cos[25007]=-78;
cos[25008]=-78;
cos[25009]=-78;
cos[25010]=-78;
cos[25011]=-78;
cos[25012]=-78;
cos[25013]=-78;
cos[25014]=-78;
cos[25015]=-78;
cos[25016]=-78;
cos[25017]=-78;
cos[25018]=-78;
cos[25019]=-78;
cos[25020]=-78;
cos[25021]=-78;
cos[25022]=-78;
cos[25023]=-78;
cos[25024]=-78;
cos[25025]=-78;
cos[25026]=-78;
cos[25027]=-78;
cos[25028]=-78;
cos[25029]=-78;
cos[25030]=-78;
cos[25031]=-78;
cos[25032]=-78;
cos[25033]=-78;
cos[25034]=-78;
cos[25035]=-78;
cos[25036]=-78;
cos[25037]=-78;
cos[25038]=-78;
cos[25039]=-78;
cos[25040]=-78;
cos[25041]=-78;
cos[25042]=-78;
cos[25043]=-78;
cos[25044]=-78;
cos[25045]=-78;
cos[25046]=-78;
cos[25047]=-78;
cos[25048]=-78;
cos[25049]=-78;
cos[25050]=-78;
cos[25051]=-78;
cos[25052]=-78;
cos[25053]=-78;
cos[25054]=-78;
cos[25055]=-78;
cos[25056]=-78;
cos[25057]=-78;
cos[25058]=-78;
cos[25059]=-78;
cos[25060]=-78;
cos[25061]=-78;
cos[25062]=-78;
cos[25063]=-78;
cos[25064]=-78;
cos[25065]=-78;
cos[25066]=-78;
cos[25067]=-78;
cos[25068]=-78;
cos[25069]=-78;
cos[25070]=-78;
cos[25071]=-78;
cos[25072]=-78;
cos[25073]=-78;
cos[25074]=-78;
cos[25075]=-78;
cos[25076]=-78;
cos[25077]=-78;
cos[25078]=-78;
cos[25079]=-78;
cos[25080]=-78;
cos[25081]=-78;
cos[25082]=-78;
cos[25083]=-78;
cos[25084]=-78;
cos[25085]=-78;
cos[25086]=-78;
cos[25087]=-78;
cos[25088]=-78;
cos[25089]=-78;
cos[25090]=-78;
cos[25091]=-78;
cos[25092]=-78;
cos[25093]=-78;
cos[25094]=-78;
cos[25095]=-78;
cos[25096]=-78;
cos[25097]=-78;
cos[25098]=-78;
cos[25099]=-78;
cos[25100]=-78;
cos[25101]=-78;
cos[25102]=-78;
cos[25103]=-78;
cos[25104]=-78;
cos[25105]=-78;
cos[25106]=-78;
cos[25107]=-78;
cos[25108]=-78;
cos[25109]=-78;
cos[25110]=-78;
cos[25111]=-78;
cos[25112]=-78;
cos[25113]=-78;
cos[25114]=-78;
cos[25115]=-78;
cos[25116]=-78;
cos[25117]=-78;
cos[25118]=-78;
cos[25119]=-78;
cos[25120]=-78;
cos[25121]=-78;
cos[25122]=-78;
cos[25123]=-78;
cos[25124]=-78;
cos[25125]=-78;
cos[25126]=-78;
cos[25127]=-78;
cos[25128]=-78;
cos[25129]=-78;
cos[25130]=-78;
cos[25131]=-78;
cos[25132]=-78;
cos[25133]=-78;
cos[25134]=-78;
cos[25135]=-78;
cos[25136]=-78;
cos[25137]=-78;
cos[25138]=-78;
cos[25139]=-78;
cos[25140]=-78;
cos[25141]=-78;
cos[25142]=-78;
cos[25143]=-78;
cos[25144]=-78;
cos[25145]=-78;
cos[25146]=-78;
cos[25147]=-78;
cos[25148]=-78;
cos[25149]=-78;
cos[25150]=-78;
cos[25151]=-78;
cos[25152]=-78;
cos[25153]=-78;
cos[25154]=-78;
cos[25155]=-78;
cos[25156]=-78;
cos[25157]=-78;
cos[25158]=-78;
cos[25159]=-78;
cos[25160]=-78;
cos[25161]=-78;
cos[25162]=-78;
cos[25163]=-78;
cos[25164]=-78;
cos[25165]=-78;
cos[25166]=-78;
cos[25167]=-78;
cos[25168]=-78;
cos[25169]=-78;
cos[25170]=-78;
cos[25171]=-78;
cos[25172]=-78;
cos[25173]=-78;
cos[25174]=-78;
cos[25175]=-78;
cos[25176]=-78;
cos[25177]=-78;
cos[25178]=-78;
cos[25179]=-78;
cos[25180]=-78;
cos[25181]=-78;
cos[25182]=-78;
cos[25183]=-78;
cos[25184]=-78;
cos[25185]=-78;
cos[25186]=-78;
cos[25187]=-78;
cos[25188]=-78;
cos[25189]=-78;
cos[25190]=-78;
cos[25191]=-78;
cos[25192]=-78;
cos[25193]=-78;
cos[25194]=-78;
cos[25195]=-78;
cos[25196]=-78;
cos[25197]=-78;
cos[25198]=-78;
cos[25199]=-78;
cos[25200]=-78;
cos[25201]=-78;
cos[25202]=-77;
cos[25203]=-77;
cos[25204]=-77;
cos[25205]=-77;
cos[25206]=-77;
cos[25207]=-77;
cos[25208]=-77;
cos[25209]=-77;
cos[25210]=-77;
cos[25211]=-77;
cos[25212]=-77;
cos[25213]=-77;
cos[25214]=-77;
cos[25215]=-77;
cos[25216]=-77;
cos[25217]=-77;
cos[25218]=-77;
cos[25219]=-77;
cos[25220]=-77;
cos[25221]=-77;
cos[25222]=-77;
cos[25223]=-77;
cos[25224]=-77;
cos[25225]=-77;
cos[25226]=-77;
cos[25227]=-77;
cos[25228]=-77;
cos[25229]=-77;
cos[25230]=-77;
cos[25231]=-77;
cos[25232]=-77;
cos[25233]=-77;
cos[25234]=-77;
cos[25235]=-77;
cos[25236]=-77;
cos[25237]=-77;
cos[25238]=-77;
cos[25239]=-77;
cos[25240]=-77;
cos[25241]=-77;
cos[25242]=-77;
cos[25243]=-77;
cos[25244]=-77;
cos[25245]=-77;
cos[25246]=-77;
cos[25247]=-77;
cos[25248]=-77;
cos[25249]=-77;
cos[25250]=-77;
cos[25251]=-77;
cos[25252]=-77;
cos[25253]=-77;
cos[25254]=-77;
cos[25255]=-77;
cos[25256]=-77;
cos[25257]=-77;
cos[25258]=-77;
cos[25259]=-77;
cos[25260]=-77;
cos[25261]=-77;
cos[25262]=-77;
cos[25263]=-77;
cos[25264]=-77;
cos[25265]=-77;
cos[25266]=-77;
cos[25267]=-77;
cos[25268]=-77;
cos[25269]=-77;
cos[25270]=-77;
cos[25271]=-77;
cos[25272]=-77;
cos[25273]=-77;
cos[25274]=-77;
cos[25275]=-77;
cos[25276]=-77;
cos[25277]=-77;
cos[25278]=-77;
cos[25279]=-77;
cos[25280]=-77;
cos[25281]=-77;
cos[25282]=-77;
cos[25283]=-77;
cos[25284]=-77;
cos[25285]=-77;
cos[25286]=-77;
cos[25287]=-77;
cos[25288]=-77;
cos[25289]=-77;
cos[25290]=-77;
cos[25291]=-77;
cos[25292]=-77;
cos[25293]=-77;
cos[25294]=-77;
cos[25295]=-77;
cos[25296]=-77;
cos[25297]=-77;
cos[25298]=-77;
cos[25299]=-77;
cos[25300]=-77;
cos[25301]=-77;
cos[25302]=-77;
cos[25303]=-77;
cos[25304]=-77;
cos[25305]=-77;
cos[25306]=-77;
cos[25307]=-77;
cos[25308]=-77;
cos[25309]=-77;
cos[25310]=-77;
cos[25311]=-77;
cos[25312]=-77;
cos[25313]=-77;
cos[25314]=-77;
cos[25315]=-77;
cos[25316]=-77;
cos[25317]=-77;
cos[25318]=-77;
cos[25319]=-77;
cos[25320]=-77;
cos[25321]=-77;
cos[25322]=-77;
cos[25323]=-77;
cos[25324]=-77;
cos[25325]=-77;
cos[25326]=-76;
cos[25327]=-76;
cos[25328]=-76;
cos[25329]=-76;
cos[25330]=-76;
cos[25331]=-76;
cos[25332]=-76;
cos[25333]=-76;
cos[25334]=-76;
cos[25335]=-76;
cos[25336]=-76;
cos[25337]=-76;
cos[25338]=-76;
cos[25339]=-76;
cos[25340]=-76;
cos[25341]=-76;
cos[25342]=-76;
cos[25343]=-76;
cos[25344]=-76;
cos[25345]=-76;
cos[25346]=-76;
cos[25347]=-76;
cos[25348]=-76;
cos[25349]=-76;
cos[25350]=-76;
cos[25351]=-76;
cos[25352]=-76;
cos[25353]=-76;
cos[25354]=-76;
cos[25355]=-76;
cos[25356]=-76;
cos[25357]=-76;
cos[25358]=-76;
cos[25359]=-76;
cos[25360]=-76;
cos[25361]=-76;
cos[25362]=-76;
cos[25363]=-76;
cos[25364]=-76;
cos[25365]=-76;
cos[25366]=-76;
cos[25367]=-76;
cos[25368]=-76;
cos[25369]=-76;
cos[25370]=-76;
cos[25371]=-76;
cos[25372]=-76;
cos[25373]=-76;
cos[25374]=-76;
cos[25375]=-76;
cos[25376]=-76;
cos[25377]=-76;
cos[25378]=-76;
cos[25379]=-76;
cos[25380]=-76;
cos[25381]=-76;
cos[25382]=-76;
cos[25383]=-76;
cos[25384]=-76;
cos[25385]=-76;
cos[25386]=-76;
cos[25387]=-76;
cos[25388]=-76;
cos[25389]=-76;
cos[25390]=-76;
cos[25391]=-76;
cos[25392]=-76;
cos[25393]=-76;
cos[25394]=-76;
cos[25395]=-76;
cos[25396]=-76;
cos[25397]=-76;
cos[25398]=-76;
cos[25399]=-76;
cos[25400]=-76;
cos[25401]=-76;
cos[25402]=-76;
cos[25403]=-76;
cos[25404]=-76;
cos[25405]=-76;
cos[25406]=-76;
cos[25407]=-76;
cos[25408]=-76;
cos[25409]=-76;
cos[25410]=-76;
cos[25411]=-76;
cos[25412]=-76;
cos[25413]=-76;
cos[25414]=-75;
cos[25415]=-75;
cos[25416]=-75;
cos[25417]=-75;
cos[25418]=-75;
cos[25419]=-75;
cos[25420]=-75;
cos[25421]=-75;
cos[25422]=-75;
cos[25423]=-75;
cos[25424]=-75;
cos[25425]=-75;
cos[25426]=-75;
cos[25427]=-75;
cos[25428]=-75;
cos[25429]=-75;
cos[25430]=-75;
cos[25431]=-75;
cos[25432]=-75;
cos[25433]=-75;
cos[25434]=-75;
cos[25435]=-75;
cos[25436]=-75;
cos[25437]=-75;
cos[25438]=-75;
cos[25439]=-75;
cos[25440]=-75;
cos[25441]=-75;
cos[25442]=-75;
cos[25443]=-75;
cos[25444]=-75;
cos[25445]=-75;
cos[25446]=-75;
cos[25447]=-75;
cos[25448]=-75;
cos[25449]=-75;
cos[25450]=-75;
cos[25451]=-75;
cos[25452]=-75;
cos[25453]=-75;
cos[25454]=-75;
cos[25455]=-75;
cos[25456]=-75;
cos[25457]=-75;
cos[25458]=-75;
cos[25459]=-75;
cos[25460]=-75;
cos[25461]=-75;
cos[25462]=-75;
cos[25463]=-75;
cos[25464]=-75;
cos[25465]=-75;
cos[25466]=-75;
cos[25467]=-75;
cos[25468]=-75;
cos[25469]=-75;
cos[25470]=-75;
cos[25471]=-75;
cos[25472]=-75;
cos[25473]=-75;
cos[25474]=-75;
cos[25475]=-75;
cos[25476]=-75;
cos[25477]=-75;
cos[25478]=-75;
cos[25479]=-75;
cos[25480]=-75;
cos[25481]=-75;
cos[25482]=-75;
cos[25483]=-75;
cos[25484]=-75;
cos[25485]=-75;
cos[25486]=-75;
cos[25487]=-74;
cos[25488]=-74;
cos[25489]=-74;
cos[25490]=-74;
cos[25491]=-74;
cos[25492]=-74;
cos[25493]=-74;
cos[25494]=-74;
cos[25495]=-74;
cos[25496]=-74;
cos[25497]=-74;
cos[25498]=-74;
cos[25499]=-74;
cos[25500]=-74;
cos[25501]=-74;
cos[25502]=-74;
cos[25503]=-74;
cos[25504]=-74;
cos[25505]=-74;
cos[25506]=-74;
cos[25507]=-74;
cos[25508]=-74;
cos[25509]=-74;
cos[25510]=-74;
cos[25511]=-74;
cos[25512]=-74;
cos[25513]=-74;
cos[25514]=-74;
cos[25515]=-74;
cos[25516]=-74;
cos[25517]=-74;
cos[25518]=-74;
cos[25519]=-74;
cos[25520]=-74;
cos[25521]=-74;
cos[25522]=-74;
cos[25523]=-74;
cos[25524]=-74;
cos[25525]=-74;
cos[25526]=-74;
cos[25527]=-74;
cos[25528]=-74;
cos[25529]=-74;
cos[25530]=-74;
cos[25531]=-74;
cos[25532]=-74;
cos[25533]=-74;
cos[25534]=-74;
cos[25535]=-74;
cos[25536]=-74;
cos[25537]=-74;
cos[25538]=-74;
cos[25539]=-74;
cos[25540]=-74;
cos[25541]=-74;
cos[25542]=-74;
cos[25543]=-74;
cos[25544]=-74;
cos[25545]=-74;
cos[25546]=-74;
cos[25547]=-74;
cos[25548]=-74;
cos[25549]=-74;
cos[25550]=-74;
cos[25551]=-73;
cos[25552]=-73;
cos[25553]=-73;
cos[25554]=-73;
cos[25555]=-73;
cos[25556]=-73;
cos[25557]=-73;
cos[25558]=-73;
cos[25559]=-73;
cos[25560]=-73;
cos[25561]=-73;
cos[25562]=-73;
cos[25563]=-73;
cos[25564]=-73;
cos[25565]=-73;
cos[25566]=-73;
cos[25567]=-73;
cos[25568]=-73;
cos[25569]=-73;
cos[25570]=-73;
cos[25571]=-73;
cos[25572]=-73;
cos[25573]=-73;
cos[25574]=-73;
cos[25575]=-73;
cos[25576]=-73;
cos[25577]=-73;
cos[25578]=-73;
cos[25579]=-73;
cos[25580]=-73;
cos[25581]=-73;
cos[25582]=-73;
cos[25583]=-73;
cos[25584]=-73;
cos[25585]=-73;
cos[25586]=-73;
cos[25587]=-73;
cos[25588]=-73;
cos[25589]=-73;
cos[25590]=-73;
cos[25591]=-73;
cos[25592]=-73;
cos[25593]=-73;
cos[25594]=-73;
cos[25595]=-73;
cos[25596]=-73;
cos[25597]=-73;
cos[25598]=-73;
cos[25599]=-73;
cos[25600]=-73;
cos[25601]=-73;
cos[25602]=-73;
cos[25603]=-73;
cos[25604]=-73;
cos[25605]=-73;
cos[25606]=-73;
cos[25607]=-73;
cos[25608]=-72;
cos[25609]=-72;
cos[25610]=-72;
cos[25611]=-72;
cos[25612]=-72;
cos[25613]=-72;
cos[25614]=-72;
cos[25615]=-72;
cos[25616]=-72;
cos[25617]=-72;
cos[25618]=-72;
cos[25619]=-72;
cos[25620]=-72;
cos[25621]=-72;
cos[25622]=-72;
cos[25623]=-72;
cos[25624]=-72;
cos[25625]=-72;
cos[25626]=-72;
cos[25627]=-72;
cos[25628]=-72;
cos[25629]=-72;
cos[25630]=-72;
cos[25631]=-72;
cos[25632]=-72;
cos[25633]=-72;
cos[25634]=-72;
cos[25635]=-72;
cos[25636]=-72;
cos[25637]=-72;
cos[25638]=-72;
cos[25639]=-72;
cos[25640]=-72;
cos[25641]=-72;
cos[25642]=-72;
cos[25643]=-72;
cos[25644]=-72;
cos[25645]=-72;
cos[25646]=-72;
cos[25647]=-72;
cos[25648]=-72;
cos[25649]=-72;
cos[25650]=-72;
cos[25651]=-72;
cos[25652]=-72;
cos[25653]=-72;
cos[25654]=-72;
cos[25655]=-72;
cos[25656]=-72;
cos[25657]=-72;
cos[25658]=-72;
cos[25659]=-72;
cos[25660]=-72;
cos[25661]=-71;
cos[25662]=-71;
cos[25663]=-71;
cos[25664]=-71;
cos[25665]=-71;
cos[25666]=-71;
cos[25667]=-71;
cos[25668]=-71;
cos[25669]=-71;
cos[25670]=-71;
cos[25671]=-71;
cos[25672]=-71;
cos[25673]=-71;
cos[25674]=-71;
cos[25675]=-71;
cos[25676]=-71;
cos[25677]=-71;
cos[25678]=-71;
cos[25679]=-71;
cos[25680]=-71;
cos[25681]=-71;
cos[25682]=-71;
cos[25683]=-71;
cos[25684]=-71;
cos[25685]=-71;
cos[25686]=-71;
cos[25687]=-71;
cos[25688]=-71;
cos[25689]=-71;
cos[25690]=-71;
cos[25691]=-71;
cos[25692]=-71;
cos[25693]=-71;
cos[25694]=-71;
cos[25695]=-71;
cos[25696]=-71;
cos[25697]=-71;
cos[25698]=-71;
cos[25699]=-71;
cos[25700]=-71;
cos[25701]=-71;
cos[25702]=-71;
cos[25703]=-71;
cos[25704]=-71;
cos[25705]=-71;
cos[25706]=-71;
cos[25707]=-71;
cos[25708]=-71;
cos[25709]=-71;
cos[25710]=-70;
cos[25711]=-70;
cos[25712]=-70;
cos[25713]=-70;
cos[25714]=-70;
cos[25715]=-70;
cos[25716]=-70;
cos[25717]=-70;
cos[25718]=-70;
cos[25719]=-70;
cos[25720]=-70;
cos[25721]=-70;
cos[25722]=-70;
cos[25723]=-70;
cos[25724]=-70;
cos[25725]=-70;
cos[25726]=-70;
cos[25727]=-70;
cos[25728]=-70;
cos[25729]=-70;
cos[25730]=-70;
cos[25731]=-70;
cos[25732]=-70;
cos[25733]=-70;
cos[25734]=-70;
cos[25735]=-70;
cos[25736]=-70;
cos[25737]=-70;
cos[25738]=-70;
cos[25739]=-70;
cos[25740]=-70;
cos[25741]=-70;
cos[25742]=-70;
cos[25743]=-70;
cos[25744]=-70;
cos[25745]=-70;
cos[25746]=-70;
cos[25747]=-70;
cos[25748]=-70;
cos[25749]=-70;
cos[25750]=-70;
cos[25751]=-70;
cos[25752]=-70;
cos[25753]=-70;
cos[25754]=-70;
cos[25755]=-69;
cos[25756]=-69;
cos[25757]=-69;
cos[25758]=-69;
cos[25759]=-69;
cos[25760]=-69;
cos[25761]=-69;
cos[25762]=-69;
cos[25763]=-69;
cos[25764]=-69;
cos[25765]=-69;
cos[25766]=-69;
cos[25767]=-69;
cos[25768]=-69;
cos[25769]=-69;
cos[25770]=-69;
cos[25771]=-69;
cos[25772]=-69;
cos[25773]=-69;
cos[25774]=-69;
cos[25775]=-69;
cos[25776]=-69;
cos[25777]=-69;
cos[25778]=-69;
cos[25779]=-69;
cos[25780]=-69;
cos[25781]=-69;
cos[25782]=-69;
cos[25783]=-69;
cos[25784]=-69;
cos[25785]=-69;
cos[25786]=-69;
cos[25787]=-69;
cos[25788]=-69;
cos[25789]=-69;
cos[25790]=-69;
cos[25791]=-69;
cos[25792]=-69;
cos[25793]=-69;
cos[25794]=-69;
cos[25795]=-69;
cos[25796]=-69;
cos[25797]=-69;
cos[25798]=-69;
cos[25799]=-68;
cos[25800]=-68;
cos[25801]=-68;
cos[25802]=-68;
cos[25803]=-68;
cos[25804]=-68;
cos[25805]=-68;
cos[25806]=-68;
cos[25807]=-68;
cos[25808]=-68;
cos[25809]=-68;
cos[25810]=-68;
cos[25811]=-68;
cos[25812]=-68;
cos[25813]=-68;
cos[25814]=-68;
cos[25815]=-68;
cos[25816]=-68;
cos[25817]=-68;
cos[25818]=-68;
cos[25819]=-68;
cos[25820]=-68;
cos[25821]=-68;
cos[25822]=-68;
cos[25823]=-68;
cos[25824]=-68;
cos[25825]=-68;
cos[25826]=-68;
cos[25827]=-68;
cos[25828]=-68;
cos[25829]=-68;
cos[25830]=-68;
cos[25831]=-68;
cos[25832]=-68;
cos[25833]=-68;
cos[25834]=-68;
cos[25835]=-68;
cos[25836]=-68;
cos[25837]=-68;
cos[25838]=-68;
cos[25839]=-68;
cos[25840]=-67;
cos[25841]=-67;
cos[25842]=-67;
cos[25843]=-67;
cos[25844]=-67;
cos[25845]=-67;
cos[25846]=-67;
cos[25847]=-67;
cos[25848]=-67;
cos[25849]=-67;
cos[25850]=-67;
cos[25851]=-67;
cos[25852]=-67;
cos[25853]=-67;
cos[25854]=-67;
cos[25855]=-67;
cos[25856]=-67;
cos[25857]=-67;
cos[25858]=-67;
cos[25859]=-67;
cos[25860]=-67;
cos[25861]=-67;
cos[25862]=-67;
cos[25863]=-67;
cos[25864]=-67;
cos[25865]=-67;
cos[25866]=-67;
cos[25867]=-67;
cos[25868]=-67;
cos[25869]=-67;
cos[25870]=-67;
cos[25871]=-67;
cos[25872]=-67;
cos[25873]=-67;
cos[25874]=-67;
cos[25875]=-67;
cos[25876]=-67;
cos[25877]=-67;
cos[25878]=-67;
cos[25879]=-67;
cos[25880]=-66;
cos[25881]=-66;
cos[25882]=-66;
cos[25883]=-66;
cos[25884]=-66;
cos[25885]=-66;
cos[25886]=-66;
cos[25887]=-66;
cos[25888]=-66;
cos[25889]=-66;
cos[25890]=-66;
cos[25891]=-66;
cos[25892]=-66;
cos[25893]=-66;
cos[25894]=-66;
cos[25895]=-66;
cos[25896]=-66;
cos[25897]=-66;
cos[25898]=-66;
cos[25899]=-66;
cos[25900]=-66;
cos[25901]=-66;
cos[25902]=-66;
cos[25903]=-66;
cos[25904]=-66;
cos[25905]=-66;
cos[25906]=-66;
cos[25907]=-66;
cos[25908]=-66;
cos[25909]=-66;
cos[25910]=-66;
cos[25911]=-66;
cos[25912]=-66;
cos[25913]=-66;
cos[25914]=-66;
cos[25915]=-66;
cos[25916]=-66;
cos[25917]=-66;
cos[25918]=-65;
cos[25919]=-65;
cos[25920]=-65;
cos[25921]=-65;
cos[25922]=-65;
cos[25923]=-65;
cos[25924]=-65;
cos[25925]=-65;
cos[25926]=-65;
cos[25927]=-65;
cos[25928]=-65;
cos[25929]=-65;
cos[25930]=-65;
cos[25931]=-65;
cos[25932]=-65;
cos[25933]=-65;
cos[25934]=-65;
cos[25935]=-65;
cos[25936]=-65;
cos[25937]=-65;
cos[25938]=-65;
cos[25939]=-65;
cos[25940]=-65;
cos[25941]=-65;
cos[25942]=-65;
cos[25943]=-65;
cos[25944]=-65;
cos[25945]=-65;
cos[25946]=-65;
cos[25947]=-65;
cos[25948]=-65;
cos[25949]=-65;
cos[25950]=-65;
cos[25951]=-65;
cos[25952]=-65;
cos[25953]=-65;
cos[25954]=-65;
cos[25955]=-64;
cos[25956]=-64;
cos[25957]=-64;
cos[25958]=-64;
cos[25959]=-64;
cos[25960]=-64;
cos[25961]=-64;
cos[25962]=-64;
cos[25963]=-64;
cos[25964]=-64;
cos[25965]=-64;
cos[25966]=-64;
cos[25967]=-64;
cos[25968]=-64;
cos[25969]=-64;
cos[25970]=-64;
cos[25971]=-64;
cos[25972]=-64;
cos[25973]=-64;
cos[25974]=-64;
cos[25975]=-64;
cos[25976]=-64;
cos[25977]=-64;
cos[25978]=-64;
cos[25979]=-64;
cos[25980]=-64;
cos[25981]=-64;
cos[25982]=-64;
cos[25983]=-64;
cos[25984]=-64;
cos[25985]=-64;
cos[25986]=-64;
cos[25987]=-64;
cos[25988]=-64;
cos[25989]=-64;
cos[25990]=-63;
cos[25991]=-63;
cos[25992]=-63;
cos[25993]=-63;
cos[25994]=-63;
cos[25995]=-63;
cos[25996]=-63;
cos[25997]=-63;
cos[25998]=-63;
cos[25999]=-63;
cos[26000]=-63;
cos[26001]=-63;
cos[26002]=-63;
cos[26003]=-63;
cos[26004]=-63;
cos[26005]=-63;
cos[26006]=-63;
cos[26007]=-63;
cos[26008]=-63;
cos[26009]=-63;
cos[26010]=-63;
cos[26011]=-63;
cos[26012]=-63;
cos[26013]=-63;
cos[26014]=-63;
cos[26015]=-63;
cos[26016]=-63;
cos[26017]=-63;
cos[26018]=-63;
cos[26019]=-63;
cos[26020]=-63;
cos[26021]=-63;
cos[26022]=-63;
cos[26023]=-63;
cos[26024]=-63;
cos[26025]=-62;
cos[26026]=-62;
cos[26027]=-62;
cos[26028]=-62;
cos[26029]=-62;
cos[26030]=-62;
cos[26031]=-62;
cos[26032]=-62;
cos[26033]=-62;
cos[26034]=-62;
cos[26035]=-62;
cos[26036]=-62;
cos[26037]=-62;
cos[26038]=-62;
cos[26039]=-62;
cos[26040]=-62;
cos[26041]=-62;
cos[26042]=-62;
cos[26043]=-62;
cos[26044]=-62;
cos[26045]=-62;
cos[26046]=-62;
cos[26047]=-62;
cos[26048]=-62;
cos[26049]=-62;
cos[26050]=-62;
cos[26051]=-62;
cos[26052]=-62;
cos[26053]=-62;
cos[26054]=-62;
cos[26055]=-62;
cos[26056]=-62;
cos[26057]=-62;
cos[26058]=-61;
cos[26059]=-61;
cos[26060]=-61;
cos[26061]=-61;
cos[26062]=-61;
cos[26063]=-61;
cos[26064]=-61;
cos[26065]=-61;
cos[26066]=-61;
cos[26067]=-61;
cos[26068]=-61;
cos[26069]=-61;
cos[26070]=-61;
cos[26071]=-61;
cos[26072]=-61;
cos[26073]=-61;
cos[26074]=-61;
cos[26075]=-61;
cos[26076]=-61;
cos[26077]=-61;
cos[26078]=-61;
cos[26079]=-61;
cos[26080]=-61;
cos[26081]=-61;
cos[26082]=-61;
cos[26083]=-61;
cos[26084]=-61;
cos[26085]=-61;
cos[26086]=-61;
cos[26087]=-61;
cos[26088]=-61;
cos[26089]=-61;
cos[26090]=-61;
cos[26091]=-60;
cos[26092]=-60;
cos[26093]=-60;
cos[26094]=-60;
cos[26095]=-60;
cos[26096]=-60;
cos[26097]=-60;
cos[26098]=-60;
cos[26099]=-60;
cos[26100]=-60;
cos[26101]=-60;
cos[26102]=-60;
cos[26103]=-60;
cos[26104]=-60;
cos[26105]=-60;
cos[26106]=-60;
cos[26107]=-60;
cos[26108]=-60;
cos[26109]=-60;
cos[26110]=-60;
cos[26111]=-60;
cos[26112]=-60;
cos[26113]=-60;
cos[26114]=-60;
cos[26115]=-60;
cos[26116]=-60;
cos[26117]=-60;
cos[26118]=-60;
cos[26119]=-60;
cos[26120]=-60;
cos[26121]=-60;
cos[26122]=-60;
cos[26123]=-59;
cos[26124]=-59;
cos[26125]=-59;
cos[26126]=-59;
cos[26127]=-59;
cos[26128]=-59;
cos[26129]=-59;
cos[26130]=-59;
cos[26131]=-59;
cos[26132]=-59;
cos[26133]=-59;
cos[26134]=-59;
cos[26135]=-59;
cos[26136]=-59;
cos[26137]=-59;
cos[26138]=-59;
cos[26139]=-59;
cos[26140]=-59;
cos[26141]=-59;
cos[26142]=-59;
cos[26143]=-59;
cos[26144]=-59;
cos[26145]=-59;
cos[26146]=-59;
cos[26147]=-59;
cos[26148]=-59;
cos[26149]=-59;
cos[26150]=-59;
cos[26151]=-59;
cos[26152]=-59;
cos[26153]=-59;
cos[26154]=-58;
cos[26155]=-58;
cos[26156]=-58;
cos[26157]=-58;
cos[26158]=-58;
cos[26159]=-58;
cos[26160]=-58;
cos[26161]=-58;
cos[26162]=-58;
cos[26163]=-58;
cos[26164]=-58;
cos[26165]=-58;
cos[26166]=-58;
cos[26167]=-58;
cos[26168]=-58;
cos[26169]=-58;
cos[26170]=-58;
cos[26171]=-58;
cos[26172]=-58;
cos[26173]=-58;
cos[26174]=-58;
cos[26175]=-58;
cos[26176]=-58;
cos[26177]=-58;
cos[26178]=-58;
cos[26179]=-58;
cos[26180]=-58;
cos[26181]=-58;
cos[26182]=-58;
cos[26183]=-58;
cos[26184]=-57;
cos[26185]=-57;
cos[26186]=-57;
cos[26187]=-57;
cos[26188]=-57;
cos[26189]=-57;
cos[26190]=-57;
cos[26191]=-57;
cos[26192]=-57;
cos[26193]=-57;
cos[26194]=-57;
cos[26195]=-57;
cos[26196]=-57;
cos[26197]=-57;
cos[26198]=-57;
cos[26199]=-57;
cos[26200]=-57;
cos[26201]=-57;
cos[26202]=-57;
cos[26203]=-57;
cos[26204]=-57;
cos[26205]=-57;
cos[26206]=-57;
cos[26207]=-57;
cos[26208]=-57;
cos[26209]=-57;
cos[26210]=-57;
cos[26211]=-57;
cos[26212]=-57;
cos[26213]=-57;
cos[26214]=-56;
cos[26215]=-56;
cos[26216]=-56;
cos[26217]=-56;
cos[26218]=-56;
cos[26219]=-56;
cos[26220]=-56;
cos[26221]=-56;
cos[26222]=-56;
cos[26223]=-56;
cos[26224]=-56;
cos[26225]=-56;
cos[26226]=-56;
cos[26227]=-56;
cos[26228]=-56;
cos[26229]=-56;
cos[26230]=-56;
cos[26231]=-56;
cos[26232]=-56;
cos[26233]=-56;
cos[26234]=-56;
cos[26235]=-56;
cos[26236]=-56;
cos[26237]=-56;
cos[26238]=-56;
cos[26239]=-56;
cos[26240]=-56;
cos[26241]=-56;
cos[26242]=-56;
cos[26243]=-55;
cos[26244]=-55;
cos[26245]=-55;
cos[26246]=-55;
cos[26247]=-55;
cos[26248]=-55;
cos[26249]=-55;
cos[26250]=-55;
cos[26251]=-55;
cos[26252]=-55;
cos[26253]=-55;
cos[26254]=-55;
cos[26255]=-55;
cos[26256]=-55;
cos[26257]=-55;
cos[26258]=-55;
cos[26259]=-55;
cos[26260]=-55;
cos[26261]=-55;
cos[26262]=-55;
cos[26263]=-55;
cos[26264]=-55;
cos[26265]=-55;
cos[26266]=-55;
cos[26267]=-55;
cos[26268]=-55;
cos[26269]=-55;
cos[26270]=-55;
cos[26271]=-55;
cos[26272]=-54;
cos[26273]=-54;
cos[26274]=-54;
cos[26275]=-54;
cos[26276]=-54;
cos[26277]=-54;
cos[26278]=-54;
cos[26279]=-54;
cos[26280]=-54;
cos[26281]=-54;
cos[26282]=-54;
cos[26283]=-54;
cos[26284]=-54;
cos[26285]=-54;
cos[26286]=-54;
cos[26287]=-54;
cos[26288]=-54;
cos[26289]=-54;
cos[26290]=-54;
cos[26291]=-54;
cos[26292]=-54;
cos[26293]=-54;
cos[26294]=-54;
cos[26295]=-54;
cos[26296]=-54;
cos[26297]=-54;
cos[26298]=-54;
cos[26299]=-54;
cos[26300]=-53;
cos[26301]=-53;
cos[26302]=-53;
cos[26303]=-53;
cos[26304]=-53;
cos[26305]=-53;
cos[26306]=-53;
cos[26307]=-53;
cos[26308]=-53;
cos[26309]=-53;
cos[26310]=-53;
cos[26311]=-53;
cos[26312]=-53;
cos[26313]=-53;
cos[26314]=-53;
cos[26315]=-53;
cos[26316]=-53;
cos[26317]=-53;
cos[26318]=-53;
cos[26319]=-53;
cos[26320]=-53;
cos[26321]=-53;
cos[26322]=-53;
cos[26323]=-53;
cos[26324]=-53;
cos[26325]=-53;
cos[26326]=-53;
cos[26327]=-53;
cos[26328]=-52;
cos[26329]=-52;
cos[26330]=-52;
cos[26331]=-52;
cos[26332]=-52;
cos[26333]=-52;
cos[26334]=-52;
cos[26335]=-52;
cos[26336]=-52;
cos[26337]=-52;
cos[26338]=-52;
cos[26339]=-52;
cos[26340]=-52;
cos[26341]=-52;
cos[26342]=-52;
cos[26343]=-52;
cos[26344]=-52;
cos[26345]=-52;
cos[26346]=-52;
cos[26347]=-52;
cos[26348]=-52;
cos[26349]=-52;
cos[26350]=-52;
cos[26351]=-52;
cos[26352]=-52;
cos[26353]=-52;
cos[26354]=-52;
cos[26355]=-51;
cos[26356]=-51;
cos[26357]=-51;
cos[26358]=-51;
cos[26359]=-51;
cos[26360]=-51;
cos[26361]=-51;
cos[26362]=-51;
cos[26363]=-51;
cos[26364]=-51;
cos[26365]=-51;
cos[26366]=-51;
cos[26367]=-51;
cos[26368]=-51;
cos[26369]=-51;
cos[26370]=-51;
cos[26371]=-51;
cos[26372]=-51;
cos[26373]=-51;
cos[26374]=-51;
cos[26375]=-51;
cos[26376]=-51;
cos[26377]=-51;
cos[26378]=-51;
cos[26379]=-51;
cos[26380]=-51;
cos[26381]=-51;
cos[26382]=-50;
cos[26383]=-50;
cos[26384]=-50;
cos[26385]=-50;
cos[26386]=-50;
cos[26387]=-50;
cos[26388]=-50;
cos[26389]=-50;
cos[26390]=-50;
cos[26391]=-50;
cos[26392]=-50;
cos[26393]=-50;
cos[26394]=-50;
cos[26395]=-50;
cos[26396]=-50;
cos[26397]=-50;
cos[26398]=-50;
cos[26399]=-50;
cos[26400]=-50;
cos[26401]=-50;
cos[26402]=-50;
cos[26403]=-50;
cos[26404]=-50;
cos[26405]=-50;
cos[26406]=-50;
cos[26407]=-50;
cos[26408]=-49;
cos[26409]=-49;
cos[26410]=-49;
cos[26411]=-49;
cos[26412]=-49;
cos[26413]=-49;
cos[26414]=-49;
cos[26415]=-49;
cos[26416]=-49;
cos[26417]=-49;
cos[26418]=-49;
cos[26419]=-49;
cos[26420]=-49;
cos[26421]=-49;
cos[26422]=-49;
cos[26423]=-49;
cos[26424]=-49;
cos[26425]=-49;
cos[26426]=-49;
cos[26427]=-49;
cos[26428]=-49;
cos[26429]=-49;
cos[26430]=-49;
cos[26431]=-49;
cos[26432]=-49;
cos[26433]=-49;
cos[26434]=-49;
cos[26435]=-48;
cos[26436]=-48;
cos[26437]=-48;
cos[26438]=-48;
cos[26439]=-48;
cos[26440]=-48;
cos[26441]=-48;
cos[26442]=-48;
cos[26443]=-48;
cos[26444]=-48;
cos[26445]=-48;
cos[26446]=-48;
cos[26447]=-48;
cos[26448]=-48;
cos[26449]=-48;
cos[26450]=-48;
cos[26451]=-48;
cos[26452]=-48;
cos[26453]=-48;
cos[26454]=-48;
cos[26455]=-48;
cos[26456]=-48;
cos[26457]=-48;
cos[26458]=-48;
cos[26459]=-48;
cos[26460]=-47;
cos[26461]=-47;
cos[26462]=-47;
cos[26463]=-47;
cos[26464]=-47;
cos[26465]=-47;
cos[26466]=-47;
cos[26467]=-47;
cos[26468]=-47;
cos[26469]=-47;
cos[26470]=-47;
cos[26471]=-47;
cos[26472]=-47;
cos[26473]=-47;
cos[26474]=-47;
cos[26475]=-47;
cos[26476]=-47;
cos[26477]=-47;
cos[26478]=-47;
cos[26479]=-47;
cos[26480]=-47;
cos[26481]=-47;
cos[26482]=-47;
cos[26483]=-47;
cos[26484]=-47;
cos[26485]=-47;
cos[26486]=-46;
cos[26487]=-46;
cos[26488]=-46;
cos[26489]=-46;
cos[26490]=-46;
cos[26491]=-46;
cos[26492]=-46;
cos[26493]=-46;
cos[26494]=-46;
cos[26495]=-46;
cos[26496]=-46;
cos[26497]=-46;
cos[26498]=-46;
cos[26499]=-46;
cos[26500]=-46;
cos[26501]=-46;
cos[26502]=-46;
cos[26503]=-46;
cos[26504]=-46;
cos[26505]=-46;
cos[26506]=-46;
cos[26507]=-46;
cos[26508]=-46;
cos[26509]=-46;
cos[26510]=-46;
cos[26511]=-45;
cos[26512]=-45;
cos[26513]=-45;
cos[26514]=-45;
cos[26515]=-45;
cos[26516]=-45;
cos[26517]=-45;
cos[26518]=-45;
cos[26519]=-45;
cos[26520]=-45;
cos[26521]=-45;
cos[26522]=-45;
cos[26523]=-45;
cos[26524]=-45;
cos[26525]=-45;
cos[26526]=-45;
cos[26527]=-45;
cos[26528]=-45;
cos[26529]=-45;
cos[26530]=-45;
cos[26531]=-45;
cos[26532]=-45;
cos[26533]=-45;
cos[26534]=-45;
cos[26535]=-45;
cos[26536]=-44;
cos[26537]=-44;
cos[26538]=-44;
cos[26539]=-44;
cos[26540]=-44;
cos[26541]=-44;
cos[26542]=-44;
cos[26543]=-44;
cos[26544]=-44;
cos[26545]=-44;
cos[26546]=-44;
cos[26547]=-44;
cos[26548]=-44;
cos[26549]=-44;
cos[26550]=-44;
cos[26551]=-44;
cos[26552]=-44;
cos[26553]=-44;
cos[26554]=-44;
cos[26555]=-44;
cos[26556]=-44;
cos[26557]=-44;
cos[26558]=-44;
cos[26559]=-44;
cos[26560]=-44;
cos[26561]=-43;
cos[26562]=-43;
cos[26563]=-43;
cos[26564]=-43;
cos[26565]=-43;
cos[26566]=-43;
cos[26567]=-43;
cos[26568]=-43;
cos[26569]=-43;
cos[26570]=-43;
cos[26571]=-43;
cos[26572]=-43;
cos[26573]=-43;
cos[26574]=-43;
cos[26575]=-43;
cos[26576]=-43;
cos[26577]=-43;
cos[26578]=-43;
cos[26579]=-43;
cos[26580]=-43;
cos[26581]=-43;
cos[26582]=-43;
cos[26583]=-43;
cos[26584]=-43;
cos[26585]=-42;
cos[26586]=-42;
cos[26587]=-42;
cos[26588]=-42;
cos[26589]=-42;
cos[26590]=-42;
cos[26591]=-42;
cos[26592]=-42;
cos[26593]=-42;
cos[26594]=-42;
cos[26595]=-42;
cos[26596]=-42;
cos[26597]=-42;
cos[26598]=-42;
cos[26599]=-42;
cos[26600]=-42;
cos[26601]=-42;
cos[26602]=-42;
cos[26603]=-42;
cos[26604]=-42;
cos[26605]=-42;
cos[26606]=-42;
cos[26607]=-42;
cos[26608]=-42;
cos[26609]=-41;
cos[26610]=-41;
cos[26611]=-41;
cos[26612]=-41;
cos[26613]=-41;
cos[26614]=-41;
cos[26615]=-41;
cos[26616]=-41;
cos[26617]=-41;
cos[26618]=-41;
cos[26619]=-41;
cos[26620]=-41;
cos[26621]=-41;
cos[26622]=-41;
cos[26623]=-41;
cos[26624]=-41;
cos[26625]=-41;
cos[26626]=-41;
cos[26627]=-41;
cos[26628]=-41;
cos[26629]=-41;
cos[26630]=-41;
cos[26631]=-41;
cos[26632]=-41;
cos[26633]=-40;
cos[26634]=-40;
cos[26635]=-40;
cos[26636]=-40;
cos[26637]=-40;
cos[26638]=-40;
cos[26639]=-40;
cos[26640]=-40;
cos[26641]=-40;
cos[26642]=-40;
cos[26643]=-40;
cos[26644]=-40;
cos[26645]=-40;
cos[26646]=-40;
cos[26647]=-40;
cos[26648]=-40;
cos[26649]=-40;
cos[26650]=-40;
cos[26651]=-40;
cos[26652]=-40;
cos[26653]=-40;
cos[26654]=-40;
cos[26655]=-40;
cos[26656]=-40;
cos[26657]=-39;
cos[26658]=-39;
cos[26659]=-39;
cos[26660]=-39;
cos[26661]=-39;
cos[26662]=-39;
cos[26663]=-39;
cos[26664]=-39;
cos[26665]=-39;
cos[26666]=-39;
cos[26667]=-39;
cos[26668]=-39;
cos[26669]=-39;
cos[26670]=-39;
cos[26671]=-39;
cos[26672]=-39;
cos[26673]=-39;
cos[26674]=-39;
cos[26675]=-39;
cos[26676]=-39;
cos[26677]=-39;
cos[26678]=-39;
cos[26679]=-39;
cos[26680]=-38;
cos[26681]=-38;
cos[26682]=-38;
cos[26683]=-38;
cos[26684]=-38;
cos[26685]=-38;
cos[26686]=-38;
cos[26687]=-38;
cos[26688]=-38;
cos[26689]=-38;
cos[26690]=-38;
cos[26691]=-38;
cos[26692]=-38;
cos[26693]=-38;
cos[26694]=-38;
cos[26695]=-38;
cos[26696]=-38;
cos[26697]=-38;
cos[26698]=-38;
cos[26699]=-38;
cos[26700]=-38;
cos[26701]=-38;
cos[26702]=-38;
cos[26703]=-38;
cos[26704]=-37;
cos[26705]=-37;
cos[26706]=-37;
cos[26707]=-37;
cos[26708]=-37;
cos[26709]=-37;
cos[26710]=-37;
cos[26711]=-37;
cos[26712]=-37;
cos[26713]=-37;
cos[26714]=-37;
cos[26715]=-37;
cos[26716]=-37;
cos[26717]=-37;
cos[26718]=-37;
cos[26719]=-37;
cos[26720]=-37;
cos[26721]=-37;
cos[26722]=-37;
cos[26723]=-37;
cos[26724]=-37;
cos[26725]=-37;
cos[26726]=-37;
cos[26727]=-36;
cos[26728]=-36;
cos[26729]=-36;
cos[26730]=-36;
cos[26731]=-36;
cos[26732]=-36;
cos[26733]=-36;
cos[26734]=-36;
cos[26735]=-36;
cos[26736]=-36;
cos[26737]=-36;
cos[26738]=-36;
cos[26739]=-36;
cos[26740]=-36;
cos[26741]=-36;
cos[26742]=-36;
cos[26743]=-36;
cos[26744]=-36;
cos[26745]=-36;
cos[26746]=-36;
cos[26747]=-36;
cos[26748]=-36;
cos[26749]=-36;
cos[26750]=-35;
cos[26751]=-35;
cos[26752]=-35;
cos[26753]=-35;
cos[26754]=-35;
cos[26755]=-35;
cos[26756]=-35;
cos[26757]=-35;
cos[26758]=-35;
cos[26759]=-35;
cos[26760]=-35;
cos[26761]=-35;
cos[26762]=-35;
cos[26763]=-35;
cos[26764]=-35;
cos[26765]=-35;
cos[26766]=-35;
cos[26767]=-35;
cos[26768]=-35;
cos[26769]=-35;
cos[26770]=-35;
cos[26771]=-35;
cos[26772]=-35;
cos[26773]=-34;
cos[26774]=-34;
cos[26775]=-34;
cos[26776]=-34;
cos[26777]=-34;
cos[26778]=-34;
cos[26779]=-34;
cos[26780]=-34;
cos[26781]=-34;
cos[26782]=-34;
cos[26783]=-34;
cos[26784]=-34;
cos[26785]=-34;
cos[26786]=-34;
cos[26787]=-34;
cos[26788]=-34;
cos[26789]=-34;
cos[26790]=-34;
cos[26791]=-34;
cos[26792]=-34;
cos[26793]=-34;
cos[26794]=-34;
cos[26795]=-33;
cos[26796]=-33;
cos[26797]=-33;
cos[26798]=-33;
cos[26799]=-33;
cos[26800]=-33;
cos[26801]=-33;
cos[26802]=-33;
cos[26803]=-33;
cos[26804]=-33;
cos[26805]=-33;
cos[26806]=-33;
cos[26807]=-33;
cos[26808]=-33;
cos[26809]=-33;
cos[26810]=-33;
cos[26811]=-33;
cos[26812]=-33;
cos[26813]=-33;
cos[26814]=-33;
cos[26815]=-33;
cos[26816]=-33;
cos[26817]=-33;
cos[26818]=-32;
cos[26819]=-32;
cos[26820]=-32;
cos[26821]=-32;
cos[26822]=-32;
cos[26823]=-32;
cos[26824]=-32;
cos[26825]=-32;
cos[26826]=-32;
cos[26827]=-32;
cos[26828]=-32;
cos[26829]=-32;
cos[26830]=-32;
cos[26831]=-32;
cos[26832]=-32;
cos[26833]=-32;
cos[26834]=-32;
cos[26835]=-32;
cos[26836]=-32;
cos[26837]=-32;
cos[26838]=-32;
cos[26839]=-32;
cos[26840]=-31;
cos[26841]=-31;
cos[26842]=-31;
cos[26843]=-31;
cos[26844]=-31;
cos[26845]=-31;
cos[26846]=-31;
cos[26847]=-31;
cos[26848]=-31;
cos[26849]=-31;
cos[26850]=-31;
cos[26851]=-31;
cos[26852]=-31;
cos[26853]=-31;
cos[26854]=-31;
cos[26855]=-31;
cos[26856]=-31;
cos[26857]=-31;
cos[26858]=-31;
cos[26859]=-31;
cos[26860]=-31;
cos[26861]=-31;
cos[26862]=-30;
cos[26863]=-30;
cos[26864]=-30;
cos[26865]=-30;
cos[26866]=-30;
cos[26867]=-30;
cos[26868]=-30;
cos[26869]=-30;
cos[26870]=-30;
cos[26871]=-30;
cos[26872]=-30;
cos[26873]=-30;
cos[26874]=-30;
cos[26875]=-30;
cos[26876]=-30;
cos[26877]=-30;
cos[26878]=-30;
cos[26879]=-30;
cos[26880]=-30;
cos[26881]=-30;
cos[26882]=-30;
cos[26883]=-30;
cos[26884]=-29;
cos[26885]=-29;
cos[26886]=-29;
cos[26887]=-29;
cos[26888]=-29;
cos[26889]=-29;
cos[26890]=-29;
cos[26891]=-29;
cos[26892]=-29;
cos[26893]=-29;
cos[26894]=-29;
cos[26895]=-29;
cos[26896]=-29;
cos[26897]=-29;
cos[26898]=-29;
cos[26899]=-29;
cos[26900]=-29;
cos[26901]=-29;
cos[26902]=-29;
cos[26903]=-29;
cos[26904]=-29;
cos[26905]=-29;
cos[26906]=-28;
cos[26907]=-28;
cos[26908]=-28;
cos[26909]=-28;
cos[26910]=-28;
cos[26911]=-28;
cos[26912]=-28;
cos[26913]=-28;
cos[26914]=-28;
cos[26915]=-28;
cos[26916]=-28;
cos[26917]=-28;
cos[26918]=-28;
cos[26919]=-28;
cos[26920]=-28;
cos[26921]=-28;
cos[26922]=-28;
cos[26923]=-28;
cos[26924]=-28;
cos[26925]=-28;
cos[26926]=-28;
cos[26927]=-28;
cos[26928]=-27;
cos[26929]=-27;
cos[26930]=-27;
cos[26931]=-27;
cos[26932]=-27;
cos[26933]=-27;
cos[26934]=-27;
cos[26935]=-27;
cos[26936]=-27;
cos[26937]=-27;
cos[26938]=-27;
cos[26939]=-27;
cos[26940]=-27;
cos[26941]=-27;
cos[26942]=-27;
cos[26943]=-27;
cos[26944]=-27;
cos[26945]=-27;
cos[26946]=-27;
cos[26947]=-27;
cos[26948]=-27;
cos[26949]=-27;
cos[26950]=-26;
cos[26951]=-26;
cos[26952]=-26;
cos[26953]=-26;
cos[26954]=-26;
cos[26955]=-26;
cos[26956]=-26;
cos[26957]=-26;
cos[26958]=-26;
cos[26959]=-26;
cos[26960]=-26;
cos[26961]=-26;
cos[26962]=-26;
cos[26963]=-26;
cos[26964]=-26;
cos[26965]=-26;
cos[26966]=-26;
cos[26967]=-26;
cos[26968]=-26;
cos[26969]=-26;
cos[26970]=-26;
cos[26971]=-25;
cos[26972]=-25;
cos[26973]=-25;
cos[26974]=-25;
cos[26975]=-25;
cos[26976]=-25;
cos[26977]=-25;
cos[26978]=-25;
cos[26979]=-25;
cos[26980]=-25;
cos[26981]=-25;
cos[26982]=-25;
cos[26983]=-25;
cos[26984]=-25;
cos[26985]=-25;
cos[26986]=-25;
cos[26987]=-25;
cos[26988]=-25;
cos[26989]=-25;
cos[26990]=-25;
cos[26991]=-25;
cos[26992]=-25;
cos[26993]=-24;
cos[26994]=-24;
cos[26995]=-24;
cos[26996]=-24;
cos[26997]=-24;
cos[26998]=-24;
cos[26999]=-24;
cos[27000]=-24;
cos[27001]=-24;
cos[27002]=-24;
cos[27003]=-24;
cos[27004]=-24;
cos[27005]=-24;
cos[27006]=-24;
cos[27007]=-24;
cos[27008]=-24;
cos[27009]=-24;
cos[27010]=-24;
cos[27011]=-24;
cos[27012]=-24;
cos[27013]=-24;
cos[27014]=-23;
cos[27015]=-23;
cos[27016]=-23;
cos[27017]=-23;
cos[27018]=-23;
cos[27019]=-23;
cos[27020]=-23;
cos[27021]=-23;
cos[27022]=-23;
cos[27023]=-23;
cos[27024]=-23;
cos[27025]=-23;
cos[27026]=-23;
cos[27027]=-23;
cos[27028]=-23;
cos[27029]=-23;
cos[27030]=-23;
cos[27031]=-23;
cos[27032]=-23;
cos[27033]=-23;
cos[27034]=-23;
cos[27035]=-23;
cos[27036]=-22;
cos[27037]=-22;
cos[27038]=-22;
cos[27039]=-22;
cos[27040]=-22;
cos[27041]=-22;
cos[27042]=-22;
cos[27043]=-22;
cos[27044]=-22;
cos[27045]=-22;
cos[27046]=-22;
cos[27047]=-22;
cos[27048]=-22;
cos[27049]=-22;
cos[27050]=-22;
cos[27051]=-22;
cos[27052]=-22;
cos[27053]=-22;
cos[27054]=-22;
cos[27055]=-22;
cos[27056]=-22;
cos[27057]=-21;
cos[27058]=-21;
cos[27059]=-21;
cos[27060]=-21;
cos[27061]=-21;
cos[27062]=-21;
cos[27063]=-21;
cos[27064]=-21;
cos[27065]=-21;
cos[27066]=-21;
cos[27067]=-21;
cos[27068]=-21;
cos[27069]=-21;
cos[27070]=-21;
cos[27071]=-21;
cos[27072]=-21;
cos[27073]=-21;
cos[27074]=-21;
cos[27075]=-21;
cos[27076]=-21;
cos[27077]=-21;
cos[27078]=-20;
cos[27079]=-20;
cos[27080]=-20;
cos[27081]=-20;
cos[27082]=-20;
cos[27083]=-20;
cos[27084]=-20;
cos[27085]=-20;
cos[27086]=-20;
cos[27087]=-20;
cos[27088]=-20;
cos[27089]=-20;
cos[27090]=-20;
cos[27091]=-20;
cos[27092]=-20;
cos[27093]=-20;
cos[27094]=-20;
cos[27095]=-20;
cos[27096]=-20;
cos[27097]=-20;
cos[27098]=-20;
cos[27099]=-19;
cos[27100]=-19;
cos[27101]=-19;
cos[27102]=-19;
cos[27103]=-19;
cos[27104]=-19;
cos[27105]=-19;
cos[27106]=-19;
cos[27107]=-19;
cos[27108]=-19;
cos[27109]=-19;
cos[27110]=-19;
cos[27111]=-19;
cos[27112]=-19;
cos[27113]=-19;
cos[27114]=-19;
cos[27115]=-19;
cos[27116]=-19;
cos[27117]=-19;
cos[27118]=-19;
cos[27119]=-19;
cos[27120]=-18;
cos[27121]=-18;
cos[27122]=-18;
cos[27123]=-18;
cos[27124]=-18;
cos[27125]=-18;
cos[27126]=-18;
cos[27127]=-18;
cos[27128]=-18;
cos[27129]=-18;
cos[27130]=-18;
cos[27131]=-18;
cos[27132]=-18;
cos[27133]=-18;
cos[27134]=-18;
cos[27135]=-18;
cos[27136]=-18;
cos[27137]=-18;
cos[27138]=-18;
cos[27139]=-18;
cos[27140]=-18;
cos[27141]=-17;
cos[27142]=-17;
cos[27143]=-17;
cos[27144]=-17;
cos[27145]=-17;
cos[27146]=-17;
cos[27147]=-17;
cos[27148]=-17;
cos[27149]=-17;
cos[27150]=-17;
cos[27151]=-17;
cos[27152]=-17;
cos[27153]=-17;
cos[27154]=-17;
cos[27155]=-17;
cos[27156]=-17;
cos[27157]=-17;
cos[27158]=-17;
cos[27159]=-17;
cos[27160]=-17;
cos[27161]=-17;
cos[27162]=-16;
cos[27163]=-16;
cos[27164]=-16;
cos[27165]=-16;
cos[27166]=-16;
cos[27167]=-16;
cos[27168]=-16;
cos[27169]=-16;
cos[27170]=-16;
cos[27171]=-16;
cos[27172]=-16;
cos[27173]=-16;
cos[27174]=-16;
cos[27175]=-16;
cos[27176]=-16;
cos[27177]=-16;
cos[27178]=-16;
cos[27179]=-16;
cos[27180]=-16;
cos[27181]=-16;
cos[27182]=-16;
cos[27183]=-15;
cos[27184]=-15;
cos[27185]=-15;
cos[27186]=-15;
cos[27187]=-15;
cos[27188]=-15;
cos[27189]=-15;
cos[27190]=-15;
cos[27191]=-15;
cos[27192]=-15;
cos[27193]=-15;
cos[27194]=-15;
cos[27195]=-15;
cos[27196]=-15;
cos[27197]=-15;
cos[27198]=-15;
cos[27199]=-15;
cos[27200]=-15;
cos[27201]=-15;
cos[27202]=-15;
cos[27203]=-14;
cos[27204]=-14;
cos[27205]=-14;
cos[27206]=-14;
cos[27207]=-14;
cos[27208]=-14;
cos[27209]=-14;
cos[27210]=-14;
cos[27211]=-14;
cos[27212]=-14;
cos[27213]=-14;
cos[27214]=-14;
cos[27215]=-14;
cos[27216]=-14;
cos[27217]=-14;
cos[27218]=-14;
cos[27219]=-14;
cos[27220]=-14;
cos[27221]=-14;
cos[27222]=-14;
cos[27223]=-14;
cos[27224]=-13;
cos[27225]=-13;
cos[27226]=-13;
cos[27227]=-13;
cos[27228]=-13;
cos[27229]=-13;
cos[27230]=-13;
cos[27231]=-13;
cos[27232]=-13;
cos[27233]=-13;
cos[27234]=-13;
cos[27235]=-13;
cos[27236]=-13;
cos[27237]=-13;
cos[27238]=-13;
cos[27239]=-13;
cos[27240]=-13;
cos[27241]=-13;
cos[27242]=-13;
cos[27243]=-13;
cos[27244]=-13;
cos[27245]=-12;
cos[27246]=-12;
cos[27247]=-12;
cos[27248]=-12;
cos[27249]=-12;
cos[27250]=-12;
cos[27251]=-12;
cos[27252]=-12;
cos[27253]=-12;
cos[27254]=-12;
cos[27255]=-12;
cos[27256]=-12;
cos[27257]=-12;
cos[27258]=-12;
cos[27259]=-12;
cos[27260]=-12;
cos[27261]=-12;
cos[27262]=-12;
cos[27263]=-12;
cos[27264]=-12;
cos[27265]=-11;
cos[27266]=-11;
cos[27267]=-11;
cos[27268]=-11;
cos[27269]=-11;
cos[27270]=-11;
cos[27271]=-11;
cos[27272]=-11;
cos[27273]=-11;
cos[27274]=-11;
cos[27275]=-11;
cos[27276]=-11;
cos[27277]=-11;
cos[27278]=-11;
cos[27279]=-11;
cos[27280]=-11;
cos[27281]=-11;
cos[27282]=-11;
cos[27283]=-11;
cos[27284]=-11;
cos[27285]=-11;
cos[27286]=-10;
cos[27287]=-10;
cos[27288]=-10;
cos[27289]=-10;
cos[27290]=-10;
cos[27291]=-10;
cos[27292]=-10;
cos[27293]=-10;
cos[27294]=-10;
cos[27295]=-10;
cos[27296]=-10;
cos[27297]=-10;
cos[27298]=-10;
cos[27299]=-10;
cos[27300]=-10;
cos[27301]=-10;
cos[27302]=-10;
cos[27303]=-10;
cos[27304]=-10;
cos[27305]=-10;
cos[27306]=-9;
cos[27307]=-9;
cos[27308]=-9;
cos[27309]=-9;
cos[27310]=-9;
cos[27311]=-9;
cos[27312]=-9;
cos[27313]=-9;
cos[27314]=-9;
cos[27315]=-9;
cos[27316]=-9;
cos[27317]=-9;
cos[27318]=-9;
cos[27319]=-9;
cos[27320]=-9;
cos[27321]=-9;
cos[27322]=-9;
cos[27323]=-9;
cos[27324]=-9;
cos[27325]=-9;
cos[27326]=-9;
cos[27327]=-8;
cos[27328]=-8;
cos[27329]=-8;
cos[27330]=-8;
cos[27331]=-8;
cos[27332]=-8;
cos[27333]=-8;
cos[27334]=-8;
cos[27335]=-8;
cos[27336]=-8;
cos[27337]=-8;
cos[27338]=-8;
cos[27339]=-8;
cos[27340]=-8;
cos[27341]=-8;
cos[27342]=-8;
cos[27343]=-8;
cos[27344]=-8;
cos[27345]=-8;
cos[27346]=-8;
cos[27347]=-7;
cos[27348]=-7;
cos[27349]=-7;
cos[27350]=-7;
cos[27351]=-7;
cos[27352]=-7;
cos[27353]=-7;
cos[27354]=-7;
cos[27355]=-7;
cos[27356]=-7;
cos[27357]=-7;
cos[27358]=-7;
cos[27359]=-7;
cos[27360]=-7;
cos[27361]=-7;
cos[27362]=-7;
cos[27363]=-7;
cos[27364]=-7;
cos[27365]=-7;
cos[27366]=-7;
cos[27367]=-7;
cos[27368]=-6;
cos[27369]=-6;
cos[27370]=-6;
cos[27371]=-6;
cos[27372]=-6;
cos[27373]=-6;
cos[27374]=-6;
cos[27375]=-6;
cos[27376]=-6;
cos[27377]=-6;
cos[27378]=-6;
cos[27379]=-6;
cos[27380]=-6;
cos[27381]=-6;
cos[27382]=-6;
cos[27383]=-6;
cos[27384]=-6;
cos[27385]=-6;
cos[27386]=-6;
cos[27387]=-6;
cos[27388]=-5;
cos[27389]=-5;
cos[27390]=-5;
cos[27391]=-5;
cos[27392]=-5;
cos[27393]=-5;
cos[27394]=-5;
cos[27395]=-5;
cos[27396]=-5;
cos[27397]=-5;
cos[27398]=-5;
cos[27399]=-5;
cos[27400]=-5;
cos[27401]=-5;
cos[27402]=-5;
cos[27403]=-5;
cos[27404]=-5;
cos[27405]=-5;
cos[27406]=-5;
cos[27407]=-5;
cos[27408]=-5;
cos[27409]=-4;
cos[27410]=-4;
cos[27411]=-4;
cos[27412]=-4;
cos[27413]=-4;
cos[27414]=-4;
cos[27415]=-4;
cos[27416]=-4;
cos[27417]=-4;
cos[27418]=-4;
cos[27419]=-4;
cos[27420]=-4;
cos[27421]=-4;
cos[27422]=-4;
cos[27423]=-4;
cos[27424]=-4;
cos[27425]=-4;
cos[27426]=-4;
cos[27427]=-4;
cos[27428]=-4;
cos[27429]=-3;
cos[27430]=-3;
cos[27431]=-3;
cos[27432]=-3;
cos[27433]=-3;
cos[27434]=-3;
cos[27435]=-3;
cos[27436]=-3;
cos[27437]=-3;
cos[27438]=-3;
cos[27439]=-3;
cos[27440]=-3;
cos[27441]=-3;
cos[27442]=-3;
cos[27443]=-3;
cos[27444]=-3;
cos[27445]=-3;
cos[27446]=-3;
cos[27447]=-3;
cos[27448]=-3;
cos[27449]=-3;
cos[27450]=-2;
cos[27451]=-2;
cos[27452]=-2;
cos[27453]=-2;
cos[27454]=-2;
cos[27455]=-2;
cos[27456]=-2;
cos[27457]=-2;
cos[27458]=-2;
cos[27459]=-2;
cos[27460]=-2;
cos[27461]=-2;
cos[27462]=-2;
cos[27463]=-2;
cos[27464]=-2;
cos[27465]=-2;
cos[27466]=-2;
cos[27467]=-2;
cos[27468]=-2;
cos[27469]=-2;
cos[27470]=-1;
cos[27471]=-1;
cos[27472]=-1;
cos[27473]=-1;
cos[27474]=-1;
cos[27475]=-1;
cos[27476]=-1;
cos[27477]=-1;
cos[27478]=-1;
cos[27479]=-1;
cos[27480]=-1;
cos[27481]=-1;
cos[27482]=-1;
cos[27483]=-1;
cos[27484]=-1;
cos[27485]=-1;
cos[27486]=-1;
cos[27487]=-1;
cos[27488]=-1;
cos[27489]=-1;
cos[27490]=0;
cos[27491]=0;
cos[27492]=0;
cos[27493]=0;
cos[27494]=0;
cos[27495]=0;
cos[27496]=0;
cos[27497]=0;
cos[27498]=0;
cos[27499]=0;
cos[27500]=0;
cos[27501]=0;
cos[27502]=0;
cos[27503]=0;
cos[27504]=0;
cos[27505]=0;
cos[27506]=0;
cos[27507]=0;
cos[27508]=0;
cos[27509]=0;
cos[27510]=0;
cos[27511]=1;
cos[27512]=1;
cos[27513]=1;
cos[27514]=1;
cos[27515]=1;
cos[27516]=1;
cos[27517]=1;
cos[27518]=1;
cos[27519]=1;
cos[27520]=1;
cos[27521]=1;
cos[27522]=1;
cos[27523]=1;
cos[27524]=1;
cos[27525]=1;
cos[27526]=1;
cos[27527]=1;
cos[27528]=1;
cos[27529]=1;
cos[27530]=1;
cos[27531]=2;
cos[27532]=2;
cos[27533]=2;
cos[27534]=2;
cos[27535]=2;
cos[27536]=2;
cos[27537]=2;
cos[27538]=2;
cos[27539]=2;
cos[27540]=2;
cos[27541]=2;
cos[27542]=2;
cos[27543]=2;
cos[27544]=2;
cos[27545]=2;
cos[27546]=2;
cos[27547]=2;
cos[27548]=2;
cos[27549]=2;
cos[27550]=2;
cos[27551]=3;
cos[27552]=3;
cos[27553]=3;
cos[27554]=3;
cos[27555]=3;
cos[27556]=3;
cos[27557]=3;
cos[27558]=3;
cos[27559]=3;
cos[27560]=3;
cos[27561]=3;
cos[27562]=3;
cos[27563]=3;
cos[27564]=3;
cos[27565]=3;
cos[27566]=3;
cos[27567]=3;
cos[27568]=3;
cos[27569]=3;
cos[27570]=3;
cos[27571]=3;
cos[27572]=4;
cos[27573]=4;
cos[27574]=4;
cos[27575]=4;
cos[27576]=4;
cos[27577]=4;
cos[27578]=4;
cos[27579]=4;
cos[27580]=4;
cos[27581]=4;
cos[27582]=4;
cos[27583]=4;
cos[27584]=4;
cos[27585]=4;
cos[27586]=4;
cos[27587]=4;
cos[27588]=4;
cos[27589]=4;
cos[27590]=4;
cos[27591]=4;
cos[27592]=5;
cos[27593]=5;
cos[27594]=5;
cos[27595]=5;
cos[27596]=5;
cos[27597]=5;
cos[27598]=5;
cos[27599]=5;
cos[27600]=5;
cos[27601]=5;
cos[27602]=5;
cos[27603]=5;
cos[27604]=5;
cos[27605]=5;
cos[27606]=5;
cos[27607]=5;
cos[27608]=5;
cos[27609]=5;
cos[27610]=5;
cos[27611]=5;
cos[27612]=5;
cos[27613]=6;
cos[27614]=6;
cos[27615]=6;
cos[27616]=6;
cos[27617]=6;
cos[27618]=6;
cos[27619]=6;
cos[27620]=6;
cos[27621]=6;
cos[27622]=6;
cos[27623]=6;
cos[27624]=6;
cos[27625]=6;
cos[27626]=6;
cos[27627]=6;
cos[27628]=6;
cos[27629]=6;
cos[27630]=6;
cos[27631]=6;
cos[27632]=6;
cos[27633]=7;
cos[27634]=7;
cos[27635]=7;
cos[27636]=7;
cos[27637]=7;
cos[27638]=7;
cos[27639]=7;
cos[27640]=7;
cos[27641]=7;
cos[27642]=7;
cos[27643]=7;
cos[27644]=7;
cos[27645]=7;
cos[27646]=7;
cos[27647]=7;
cos[27648]=7;
cos[27649]=7;
cos[27650]=7;
cos[27651]=7;
cos[27652]=7;
cos[27653]=7;
cos[27654]=8;
cos[27655]=8;
cos[27656]=8;
cos[27657]=8;
cos[27658]=8;
cos[27659]=8;
cos[27660]=8;
cos[27661]=8;
cos[27662]=8;
cos[27663]=8;
cos[27664]=8;
cos[27665]=8;
cos[27666]=8;
cos[27667]=8;
cos[27668]=8;
cos[27669]=8;
cos[27670]=8;
cos[27671]=8;
cos[27672]=8;
cos[27673]=8;
cos[27674]=9;
cos[27675]=9;
cos[27676]=9;
cos[27677]=9;
cos[27678]=9;
cos[27679]=9;
cos[27680]=9;
cos[27681]=9;
cos[27682]=9;
cos[27683]=9;
cos[27684]=9;
cos[27685]=9;
cos[27686]=9;
cos[27687]=9;
cos[27688]=9;
cos[27689]=9;
cos[27690]=9;
cos[27691]=9;
cos[27692]=9;
cos[27693]=9;
cos[27694]=9;
cos[27695]=10;
cos[27696]=10;
cos[27697]=10;
cos[27698]=10;
cos[27699]=10;
cos[27700]=10;
cos[27701]=10;
cos[27702]=10;
cos[27703]=10;
cos[27704]=10;
cos[27705]=10;
cos[27706]=10;
cos[27707]=10;
cos[27708]=10;
cos[27709]=10;
cos[27710]=10;
cos[27711]=10;
cos[27712]=10;
cos[27713]=10;
cos[27714]=10;
cos[27715]=11;
cos[27716]=11;
cos[27717]=11;
cos[27718]=11;
cos[27719]=11;
cos[27720]=11;
cos[27721]=11;
cos[27722]=11;
cos[27723]=11;
cos[27724]=11;
cos[27725]=11;
cos[27726]=11;
cos[27727]=11;
cos[27728]=11;
cos[27729]=11;
cos[27730]=11;
cos[27731]=11;
cos[27732]=11;
cos[27733]=11;
cos[27734]=11;
cos[27735]=11;
cos[27736]=12;
cos[27737]=12;
cos[27738]=12;
cos[27739]=12;
cos[27740]=12;
cos[27741]=12;
cos[27742]=12;
cos[27743]=12;
cos[27744]=12;
cos[27745]=12;
cos[27746]=12;
cos[27747]=12;
cos[27748]=12;
cos[27749]=12;
cos[27750]=12;
cos[27751]=12;
cos[27752]=12;
cos[27753]=12;
cos[27754]=12;
cos[27755]=12;
cos[27756]=13;
cos[27757]=13;
cos[27758]=13;
cos[27759]=13;
cos[27760]=13;
cos[27761]=13;
cos[27762]=13;
cos[27763]=13;
cos[27764]=13;
cos[27765]=13;
cos[27766]=13;
cos[27767]=13;
cos[27768]=13;
cos[27769]=13;
cos[27770]=13;
cos[27771]=13;
cos[27772]=13;
cos[27773]=13;
cos[27774]=13;
cos[27775]=13;
cos[27776]=13;
cos[27777]=14;
cos[27778]=14;
cos[27779]=14;
cos[27780]=14;
cos[27781]=14;
cos[27782]=14;
cos[27783]=14;
cos[27784]=14;
cos[27785]=14;
cos[27786]=14;
cos[27787]=14;
cos[27788]=14;
cos[27789]=14;
cos[27790]=14;
cos[27791]=14;
cos[27792]=14;
cos[27793]=14;
cos[27794]=14;
cos[27795]=14;
cos[27796]=14;
cos[27797]=14;
cos[27798]=15;
cos[27799]=15;
cos[27800]=15;
cos[27801]=15;
cos[27802]=15;
cos[27803]=15;
cos[27804]=15;
cos[27805]=15;
cos[27806]=15;
cos[27807]=15;
cos[27808]=15;
cos[27809]=15;
cos[27810]=15;
cos[27811]=15;
cos[27812]=15;
cos[27813]=15;
cos[27814]=15;
cos[27815]=15;
cos[27816]=15;
cos[27817]=15;
cos[27818]=16;
cos[27819]=16;
cos[27820]=16;
cos[27821]=16;
cos[27822]=16;
cos[27823]=16;
cos[27824]=16;
cos[27825]=16;
cos[27826]=16;
cos[27827]=16;
cos[27828]=16;
cos[27829]=16;
cos[27830]=16;
cos[27831]=16;
cos[27832]=16;
cos[27833]=16;
cos[27834]=16;
cos[27835]=16;
cos[27836]=16;
cos[27837]=16;
cos[27838]=16;
cos[27839]=17;
cos[27840]=17;
cos[27841]=17;
cos[27842]=17;
cos[27843]=17;
cos[27844]=17;
cos[27845]=17;
cos[27846]=17;
cos[27847]=17;
cos[27848]=17;
cos[27849]=17;
cos[27850]=17;
cos[27851]=17;
cos[27852]=17;
cos[27853]=17;
cos[27854]=17;
cos[27855]=17;
cos[27856]=17;
cos[27857]=17;
cos[27858]=17;
cos[27859]=17;
cos[27860]=18;
cos[27861]=18;
cos[27862]=18;
cos[27863]=18;
cos[27864]=18;
cos[27865]=18;
cos[27866]=18;
cos[27867]=18;
cos[27868]=18;
cos[27869]=18;
cos[27870]=18;
cos[27871]=18;
cos[27872]=18;
cos[27873]=18;
cos[27874]=18;
cos[27875]=18;
cos[27876]=18;
cos[27877]=18;
cos[27878]=18;
cos[27879]=18;
cos[27880]=18;
cos[27881]=19;
cos[27882]=19;
cos[27883]=19;
cos[27884]=19;
cos[27885]=19;
cos[27886]=19;
cos[27887]=19;
cos[27888]=19;
cos[27889]=19;
cos[27890]=19;
cos[27891]=19;
cos[27892]=19;
cos[27893]=19;
cos[27894]=19;
cos[27895]=19;
cos[27896]=19;
cos[27897]=19;
cos[27898]=19;
cos[27899]=19;
cos[27900]=19;
cos[27901]=19;
cos[27902]=20;
cos[27903]=20;
cos[27904]=20;
cos[27905]=20;
cos[27906]=20;
cos[27907]=20;
cos[27908]=20;
cos[27909]=20;
cos[27910]=20;
cos[27911]=20;
cos[27912]=20;
cos[27913]=20;
cos[27914]=20;
cos[27915]=20;
cos[27916]=20;
cos[27917]=20;
cos[27918]=20;
cos[27919]=20;
cos[27920]=20;
cos[27921]=20;
cos[27922]=20;
cos[27923]=21;
cos[27924]=21;
cos[27925]=21;
cos[27926]=21;
cos[27927]=21;
cos[27928]=21;
cos[27929]=21;
cos[27930]=21;
cos[27931]=21;
cos[27932]=21;
cos[27933]=21;
cos[27934]=21;
cos[27935]=21;
cos[27936]=21;
cos[27937]=21;
cos[27938]=21;
cos[27939]=21;
cos[27940]=21;
cos[27941]=21;
cos[27942]=21;
cos[27943]=21;
cos[27944]=22;
cos[27945]=22;
cos[27946]=22;
cos[27947]=22;
cos[27948]=22;
cos[27949]=22;
cos[27950]=22;
cos[27951]=22;
cos[27952]=22;
cos[27953]=22;
cos[27954]=22;
cos[27955]=22;
cos[27956]=22;
cos[27957]=22;
cos[27958]=22;
cos[27959]=22;
cos[27960]=22;
cos[27961]=22;
cos[27962]=22;
cos[27963]=22;
cos[27964]=22;
cos[27965]=23;
cos[27966]=23;
cos[27967]=23;
cos[27968]=23;
cos[27969]=23;
cos[27970]=23;
cos[27971]=23;
cos[27972]=23;
cos[27973]=23;
cos[27974]=23;
cos[27975]=23;
cos[27976]=23;
cos[27977]=23;
cos[27978]=23;
cos[27979]=23;
cos[27980]=23;
cos[27981]=23;
cos[27982]=23;
cos[27983]=23;
cos[27984]=23;
cos[27985]=23;
cos[27986]=23;
cos[27987]=24;
cos[27988]=24;
cos[27989]=24;
cos[27990]=24;
cos[27991]=24;
cos[27992]=24;
cos[27993]=24;
cos[27994]=24;
cos[27995]=24;
cos[27996]=24;
cos[27997]=24;
cos[27998]=24;
cos[27999]=24;
cos[28000]=24;
cos[28001]=24;
cos[28002]=24;
cos[28003]=24;
cos[28004]=24;
cos[28005]=24;
cos[28006]=24;
cos[28007]=24;
cos[28008]=25;
cos[28009]=25;
cos[28010]=25;
cos[28011]=25;
cos[28012]=25;
cos[28013]=25;
cos[28014]=25;
cos[28015]=25;
cos[28016]=25;
cos[28017]=25;
cos[28018]=25;
cos[28019]=25;
cos[28020]=25;
cos[28021]=25;
cos[28022]=25;
cos[28023]=25;
cos[28024]=25;
cos[28025]=25;
cos[28026]=25;
cos[28027]=25;
cos[28028]=25;
cos[28029]=25;
cos[28030]=26;
cos[28031]=26;
cos[28032]=26;
cos[28033]=26;
cos[28034]=26;
cos[28035]=26;
cos[28036]=26;
cos[28037]=26;
cos[28038]=26;
cos[28039]=26;
cos[28040]=26;
cos[28041]=26;
cos[28042]=26;
cos[28043]=26;
cos[28044]=26;
cos[28045]=26;
cos[28046]=26;
cos[28047]=26;
cos[28048]=26;
cos[28049]=26;
cos[28050]=26;
cos[28051]=27;
cos[28052]=27;
cos[28053]=27;
cos[28054]=27;
cos[28055]=27;
cos[28056]=27;
cos[28057]=27;
cos[28058]=27;
cos[28059]=27;
cos[28060]=27;
cos[28061]=27;
cos[28062]=27;
cos[28063]=27;
cos[28064]=27;
cos[28065]=27;
cos[28066]=27;
cos[28067]=27;
cos[28068]=27;
cos[28069]=27;
cos[28070]=27;
cos[28071]=27;
cos[28072]=27;
cos[28073]=28;
cos[28074]=28;
cos[28075]=28;
cos[28076]=28;
cos[28077]=28;
cos[28078]=28;
cos[28079]=28;
cos[28080]=28;
cos[28081]=28;
cos[28082]=28;
cos[28083]=28;
cos[28084]=28;
cos[28085]=28;
cos[28086]=28;
cos[28087]=28;
cos[28088]=28;
cos[28089]=28;
cos[28090]=28;
cos[28091]=28;
cos[28092]=28;
cos[28093]=28;
cos[28094]=28;
cos[28095]=29;
cos[28096]=29;
cos[28097]=29;
cos[28098]=29;
cos[28099]=29;
cos[28100]=29;
cos[28101]=29;
cos[28102]=29;
cos[28103]=29;
cos[28104]=29;
cos[28105]=29;
cos[28106]=29;
cos[28107]=29;
cos[28108]=29;
cos[28109]=29;
cos[28110]=29;
cos[28111]=29;
cos[28112]=29;
cos[28113]=29;
cos[28114]=29;
cos[28115]=29;
cos[28116]=29;
cos[28117]=30;
cos[28118]=30;
cos[28119]=30;
cos[28120]=30;
cos[28121]=30;
cos[28122]=30;
cos[28123]=30;
cos[28124]=30;
cos[28125]=30;
cos[28126]=30;
cos[28127]=30;
cos[28128]=30;
cos[28129]=30;
cos[28130]=30;
cos[28131]=30;
cos[28132]=30;
cos[28133]=30;
cos[28134]=30;
cos[28135]=30;
cos[28136]=30;
cos[28137]=30;
cos[28138]=30;
cos[28139]=31;
cos[28140]=31;
cos[28141]=31;
cos[28142]=31;
cos[28143]=31;
cos[28144]=31;
cos[28145]=31;
cos[28146]=31;
cos[28147]=31;
cos[28148]=31;
cos[28149]=31;
cos[28150]=31;
cos[28151]=31;
cos[28152]=31;
cos[28153]=31;
cos[28154]=31;
cos[28155]=31;
cos[28156]=31;
cos[28157]=31;
cos[28158]=31;
cos[28159]=31;
cos[28160]=31;
cos[28161]=32;
cos[28162]=32;
cos[28163]=32;
cos[28164]=32;
cos[28165]=32;
cos[28166]=32;
cos[28167]=32;
cos[28168]=32;
cos[28169]=32;
cos[28170]=32;
cos[28171]=32;
cos[28172]=32;
cos[28173]=32;
cos[28174]=32;
cos[28175]=32;
cos[28176]=32;
cos[28177]=32;
cos[28178]=32;
cos[28179]=32;
cos[28180]=32;
cos[28181]=32;
cos[28182]=32;
cos[28183]=33;
cos[28184]=33;
cos[28185]=33;
cos[28186]=33;
cos[28187]=33;
cos[28188]=33;
cos[28189]=33;
cos[28190]=33;
cos[28191]=33;
cos[28192]=33;
cos[28193]=33;
cos[28194]=33;
cos[28195]=33;
cos[28196]=33;
cos[28197]=33;
cos[28198]=33;
cos[28199]=33;
cos[28200]=33;
cos[28201]=33;
cos[28202]=33;
cos[28203]=33;
cos[28204]=33;
cos[28205]=33;
cos[28206]=34;
cos[28207]=34;
cos[28208]=34;
cos[28209]=34;
cos[28210]=34;
cos[28211]=34;
cos[28212]=34;
cos[28213]=34;
cos[28214]=34;
cos[28215]=34;
cos[28216]=34;
cos[28217]=34;
cos[28218]=34;
cos[28219]=34;
cos[28220]=34;
cos[28221]=34;
cos[28222]=34;
cos[28223]=34;
cos[28224]=34;
cos[28225]=34;
cos[28226]=34;
cos[28227]=34;
cos[28228]=35;
cos[28229]=35;
cos[28230]=35;
cos[28231]=35;
cos[28232]=35;
cos[28233]=35;
cos[28234]=35;
cos[28235]=35;
cos[28236]=35;
cos[28237]=35;
cos[28238]=35;
cos[28239]=35;
cos[28240]=35;
cos[28241]=35;
cos[28242]=35;
cos[28243]=35;
cos[28244]=35;
cos[28245]=35;
cos[28246]=35;
cos[28247]=35;
cos[28248]=35;
cos[28249]=35;
cos[28250]=35;
cos[28251]=36;
cos[28252]=36;
cos[28253]=36;
cos[28254]=36;
cos[28255]=36;
cos[28256]=36;
cos[28257]=36;
cos[28258]=36;
cos[28259]=36;
cos[28260]=36;
cos[28261]=36;
cos[28262]=36;
cos[28263]=36;
cos[28264]=36;
cos[28265]=36;
cos[28266]=36;
cos[28267]=36;
cos[28268]=36;
cos[28269]=36;
cos[28270]=36;
cos[28271]=36;
cos[28272]=36;
cos[28273]=36;
cos[28274]=37;
cos[28275]=37;
cos[28276]=37;
cos[28277]=37;
cos[28278]=37;
cos[28279]=37;
cos[28280]=37;
cos[28281]=37;
cos[28282]=37;
cos[28283]=37;
cos[28284]=37;
cos[28285]=37;
cos[28286]=37;
cos[28287]=37;
cos[28288]=37;
cos[28289]=37;
cos[28290]=37;
cos[28291]=37;
cos[28292]=37;
cos[28293]=37;
cos[28294]=37;
cos[28295]=37;
cos[28296]=37;
cos[28297]=38;
cos[28298]=38;
cos[28299]=38;
cos[28300]=38;
cos[28301]=38;
cos[28302]=38;
cos[28303]=38;
cos[28304]=38;
cos[28305]=38;
cos[28306]=38;
cos[28307]=38;
cos[28308]=38;
cos[28309]=38;
cos[28310]=38;
cos[28311]=38;
cos[28312]=38;
cos[28313]=38;
cos[28314]=38;
cos[28315]=38;
cos[28316]=38;
cos[28317]=38;
cos[28318]=38;
cos[28319]=38;
cos[28320]=38;
cos[28321]=39;
cos[28322]=39;
cos[28323]=39;
cos[28324]=39;
cos[28325]=39;
cos[28326]=39;
cos[28327]=39;
cos[28328]=39;
cos[28329]=39;
cos[28330]=39;
cos[28331]=39;
cos[28332]=39;
cos[28333]=39;
cos[28334]=39;
cos[28335]=39;
cos[28336]=39;
cos[28337]=39;
cos[28338]=39;
cos[28339]=39;
cos[28340]=39;
cos[28341]=39;
cos[28342]=39;
cos[28343]=39;
cos[28344]=40;
cos[28345]=40;
cos[28346]=40;
cos[28347]=40;
cos[28348]=40;
cos[28349]=40;
cos[28350]=40;
cos[28351]=40;
cos[28352]=40;
cos[28353]=40;
cos[28354]=40;
cos[28355]=40;
cos[28356]=40;
cos[28357]=40;
cos[28358]=40;
cos[28359]=40;
cos[28360]=40;
cos[28361]=40;
cos[28362]=40;
cos[28363]=40;
cos[28364]=40;
cos[28365]=40;
cos[28366]=40;
cos[28367]=40;
cos[28368]=41;
cos[28369]=41;
cos[28370]=41;
cos[28371]=41;
cos[28372]=41;
cos[28373]=41;
cos[28374]=41;
cos[28375]=41;
cos[28376]=41;
cos[28377]=41;
cos[28378]=41;
cos[28379]=41;
cos[28380]=41;
cos[28381]=41;
cos[28382]=41;
cos[28383]=41;
cos[28384]=41;
cos[28385]=41;
cos[28386]=41;
cos[28387]=41;
cos[28388]=41;
cos[28389]=41;
cos[28390]=41;
cos[28391]=41;
cos[28392]=42;
cos[28393]=42;
cos[28394]=42;
cos[28395]=42;
cos[28396]=42;
cos[28397]=42;
cos[28398]=42;
cos[28399]=42;
cos[28400]=42;
cos[28401]=42;
cos[28402]=42;
cos[28403]=42;
cos[28404]=42;
cos[28405]=42;
cos[28406]=42;
cos[28407]=42;
cos[28408]=42;
cos[28409]=42;
cos[28410]=42;
cos[28411]=42;
cos[28412]=42;
cos[28413]=42;
cos[28414]=42;
cos[28415]=42;
cos[28416]=43;
cos[28417]=43;
cos[28418]=43;
cos[28419]=43;
cos[28420]=43;
cos[28421]=43;
cos[28422]=43;
cos[28423]=43;
cos[28424]=43;
cos[28425]=43;
cos[28426]=43;
cos[28427]=43;
cos[28428]=43;
cos[28429]=43;
cos[28430]=43;
cos[28431]=43;
cos[28432]=43;
cos[28433]=43;
cos[28434]=43;
cos[28435]=43;
cos[28436]=43;
cos[28437]=43;
cos[28438]=43;
cos[28439]=43;
cos[28440]=44;
cos[28441]=44;
cos[28442]=44;
cos[28443]=44;
cos[28444]=44;
cos[28445]=44;
cos[28446]=44;
cos[28447]=44;
cos[28448]=44;
cos[28449]=44;
cos[28450]=44;
cos[28451]=44;
cos[28452]=44;
cos[28453]=44;
cos[28454]=44;
cos[28455]=44;
cos[28456]=44;
cos[28457]=44;
cos[28458]=44;
cos[28459]=44;
cos[28460]=44;
cos[28461]=44;
cos[28462]=44;
cos[28463]=44;
cos[28464]=44;
cos[28465]=45;
cos[28466]=45;
cos[28467]=45;
cos[28468]=45;
cos[28469]=45;
cos[28470]=45;
cos[28471]=45;
cos[28472]=45;
cos[28473]=45;
cos[28474]=45;
cos[28475]=45;
cos[28476]=45;
cos[28477]=45;
cos[28478]=45;
cos[28479]=45;
cos[28480]=45;
cos[28481]=45;
cos[28482]=45;
cos[28483]=45;
cos[28484]=45;
cos[28485]=45;
cos[28486]=45;
cos[28487]=45;
cos[28488]=45;
cos[28489]=45;
cos[28490]=46;
cos[28491]=46;
cos[28492]=46;
cos[28493]=46;
cos[28494]=46;
cos[28495]=46;
cos[28496]=46;
cos[28497]=46;
cos[28498]=46;
cos[28499]=46;
cos[28500]=46;
cos[28501]=46;
cos[28502]=46;
cos[28503]=46;
cos[28504]=46;
cos[28505]=46;
cos[28506]=46;
cos[28507]=46;
cos[28508]=46;
cos[28509]=46;
cos[28510]=46;
cos[28511]=46;
cos[28512]=46;
cos[28513]=46;
cos[28514]=46;
cos[28515]=47;
cos[28516]=47;
cos[28517]=47;
cos[28518]=47;
cos[28519]=47;
cos[28520]=47;
cos[28521]=47;
cos[28522]=47;
cos[28523]=47;
cos[28524]=47;
cos[28525]=47;
cos[28526]=47;
cos[28527]=47;
cos[28528]=47;
cos[28529]=47;
cos[28530]=47;
cos[28531]=47;
cos[28532]=47;
cos[28533]=47;
cos[28534]=47;
cos[28535]=47;
cos[28536]=47;
cos[28537]=47;
cos[28538]=47;
cos[28539]=47;
cos[28540]=47;
cos[28541]=48;
cos[28542]=48;
cos[28543]=48;
cos[28544]=48;
cos[28545]=48;
cos[28546]=48;
cos[28547]=48;
cos[28548]=48;
cos[28549]=48;
cos[28550]=48;
cos[28551]=48;
cos[28552]=48;
cos[28553]=48;
cos[28554]=48;
cos[28555]=48;
cos[28556]=48;
cos[28557]=48;
cos[28558]=48;
cos[28559]=48;
cos[28560]=48;
cos[28561]=48;
cos[28562]=48;
cos[28563]=48;
cos[28564]=48;
cos[28565]=48;
cos[28566]=49;
cos[28567]=49;
cos[28568]=49;
cos[28569]=49;
cos[28570]=49;
cos[28571]=49;
cos[28572]=49;
cos[28573]=49;
cos[28574]=49;
cos[28575]=49;
cos[28576]=49;
cos[28577]=49;
cos[28578]=49;
cos[28579]=49;
cos[28580]=49;
cos[28581]=49;
cos[28582]=49;
cos[28583]=49;
cos[28584]=49;
cos[28585]=49;
cos[28586]=49;
cos[28587]=49;
cos[28588]=49;
cos[28589]=49;
cos[28590]=49;
cos[28591]=49;
cos[28592]=49;
cos[28593]=50;
cos[28594]=50;
cos[28595]=50;
cos[28596]=50;
cos[28597]=50;
cos[28598]=50;
cos[28599]=50;
cos[28600]=50;
cos[28601]=50;
cos[28602]=50;
cos[28603]=50;
cos[28604]=50;
cos[28605]=50;
cos[28606]=50;
cos[28607]=50;
cos[28608]=50;
cos[28609]=50;
cos[28610]=50;
cos[28611]=50;
cos[28612]=50;
cos[28613]=50;
cos[28614]=50;
cos[28615]=50;
cos[28616]=50;
cos[28617]=50;
cos[28618]=50;
cos[28619]=51;
cos[28620]=51;
cos[28621]=51;
cos[28622]=51;
cos[28623]=51;
cos[28624]=51;
cos[28625]=51;
cos[28626]=51;
cos[28627]=51;
cos[28628]=51;
cos[28629]=51;
cos[28630]=51;
cos[28631]=51;
cos[28632]=51;
cos[28633]=51;
cos[28634]=51;
cos[28635]=51;
cos[28636]=51;
cos[28637]=51;
cos[28638]=51;
cos[28639]=51;
cos[28640]=51;
cos[28641]=51;
cos[28642]=51;
cos[28643]=51;
cos[28644]=51;
cos[28645]=51;
cos[28646]=52;
cos[28647]=52;
cos[28648]=52;
cos[28649]=52;
cos[28650]=52;
cos[28651]=52;
cos[28652]=52;
cos[28653]=52;
cos[28654]=52;
cos[28655]=52;
cos[28656]=52;
cos[28657]=52;
cos[28658]=52;
cos[28659]=52;
cos[28660]=52;
cos[28661]=52;
cos[28662]=52;
cos[28663]=52;
cos[28664]=52;
cos[28665]=52;
cos[28666]=52;
cos[28667]=52;
cos[28668]=52;
cos[28669]=52;
cos[28670]=52;
cos[28671]=52;
cos[28672]=52;
cos[28673]=53;
cos[28674]=53;
cos[28675]=53;
cos[28676]=53;
cos[28677]=53;
cos[28678]=53;
cos[28679]=53;
cos[28680]=53;
cos[28681]=53;
cos[28682]=53;
cos[28683]=53;
cos[28684]=53;
cos[28685]=53;
cos[28686]=53;
cos[28687]=53;
cos[28688]=53;
cos[28689]=53;
cos[28690]=53;
cos[28691]=53;
cos[28692]=53;
cos[28693]=53;
cos[28694]=53;
cos[28695]=53;
cos[28696]=53;
cos[28697]=53;
cos[28698]=53;
cos[28699]=53;
cos[28700]=53;
cos[28701]=54;
cos[28702]=54;
cos[28703]=54;
cos[28704]=54;
cos[28705]=54;
cos[28706]=54;
cos[28707]=54;
cos[28708]=54;
cos[28709]=54;
cos[28710]=54;
cos[28711]=54;
cos[28712]=54;
cos[28713]=54;
cos[28714]=54;
cos[28715]=54;
cos[28716]=54;
cos[28717]=54;
cos[28718]=54;
cos[28719]=54;
cos[28720]=54;
cos[28721]=54;
cos[28722]=54;
cos[28723]=54;
cos[28724]=54;
cos[28725]=54;
cos[28726]=54;
cos[28727]=54;
cos[28728]=54;
cos[28729]=55;
cos[28730]=55;
cos[28731]=55;
cos[28732]=55;
cos[28733]=55;
cos[28734]=55;
cos[28735]=55;
cos[28736]=55;
cos[28737]=55;
cos[28738]=55;
cos[28739]=55;
cos[28740]=55;
cos[28741]=55;
cos[28742]=55;
cos[28743]=55;
cos[28744]=55;
cos[28745]=55;
cos[28746]=55;
cos[28747]=55;
cos[28748]=55;
cos[28749]=55;
cos[28750]=55;
cos[28751]=55;
cos[28752]=55;
cos[28753]=55;
cos[28754]=55;
cos[28755]=55;
cos[28756]=55;
cos[28757]=55;
cos[28758]=56;
cos[28759]=56;
cos[28760]=56;
cos[28761]=56;
cos[28762]=56;
cos[28763]=56;
cos[28764]=56;
cos[28765]=56;
cos[28766]=56;
cos[28767]=56;
cos[28768]=56;
cos[28769]=56;
cos[28770]=56;
cos[28771]=56;
cos[28772]=56;
cos[28773]=56;
cos[28774]=56;
cos[28775]=56;
cos[28776]=56;
cos[28777]=56;
cos[28778]=56;
cos[28779]=56;
cos[28780]=56;
cos[28781]=56;
cos[28782]=56;
cos[28783]=56;
cos[28784]=56;
cos[28785]=56;
cos[28786]=56;
cos[28787]=57;
cos[28788]=57;
cos[28789]=57;
cos[28790]=57;
cos[28791]=57;
cos[28792]=57;
cos[28793]=57;
cos[28794]=57;
cos[28795]=57;
cos[28796]=57;
cos[28797]=57;
cos[28798]=57;
cos[28799]=57;
cos[28800]=57;
cos[28801]=57;
cos[28802]=57;
cos[28803]=57;
cos[28804]=57;
cos[28805]=57;
cos[28806]=57;
cos[28807]=57;
cos[28808]=57;
cos[28809]=57;
cos[28810]=57;
cos[28811]=57;
cos[28812]=57;
cos[28813]=57;
cos[28814]=57;
cos[28815]=57;
cos[28816]=57;
cos[28817]=58;
cos[28818]=58;
cos[28819]=58;
cos[28820]=58;
cos[28821]=58;
cos[28822]=58;
cos[28823]=58;
cos[28824]=58;
cos[28825]=58;
cos[28826]=58;
cos[28827]=58;
cos[28828]=58;
cos[28829]=58;
cos[28830]=58;
cos[28831]=58;
cos[28832]=58;
cos[28833]=58;
cos[28834]=58;
cos[28835]=58;
cos[28836]=58;
cos[28837]=58;
cos[28838]=58;
cos[28839]=58;
cos[28840]=58;
cos[28841]=58;
cos[28842]=58;
cos[28843]=58;
cos[28844]=58;
cos[28845]=58;
cos[28846]=58;
cos[28847]=59;
cos[28848]=59;
cos[28849]=59;
cos[28850]=59;
cos[28851]=59;
cos[28852]=59;
cos[28853]=59;
cos[28854]=59;
cos[28855]=59;
cos[28856]=59;
cos[28857]=59;
cos[28858]=59;
cos[28859]=59;
cos[28860]=59;
cos[28861]=59;
cos[28862]=59;
cos[28863]=59;
cos[28864]=59;
cos[28865]=59;
cos[28866]=59;
cos[28867]=59;
cos[28868]=59;
cos[28869]=59;
cos[28870]=59;
cos[28871]=59;
cos[28872]=59;
cos[28873]=59;
cos[28874]=59;
cos[28875]=59;
cos[28876]=59;
cos[28877]=59;
cos[28878]=60;
cos[28879]=60;
cos[28880]=60;
cos[28881]=60;
cos[28882]=60;
cos[28883]=60;
cos[28884]=60;
cos[28885]=60;
cos[28886]=60;
cos[28887]=60;
cos[28888]=60;
cos[28889]=60;
cos[28890]=60;
cos[28891]=60;
cos[28892]=60;
cos[28893]=60;
cos[28894]=60;
cos[28895]=60;
cos[28896]=60;
cos[28897]=60;
cos[28898]=60;
cos[28899]=60;
cos[28900]=60;
cos[28901]=60;
cos[28902]=60;
cos[28903]=60;
cos[28904]=60;
cos[28905]=60;
cos[28906]=60;
cos[28907]=60;
cos[28908]=60;
cos[28909]=60;
cos[28910]=61;
cos[28911]=61;
cos[28912]=61;
cos[28913]=61;
cos[28914]=61;
cos[28915]=61;
cos[28916]=61;
cos[28917]=61;
cos[28918]=61;
cos[28919]=61;
cos[28920]=61;
cos[28921]=61;
cos[28922]=61;
cos[28923]=61;
cos[28924]=61;
cos[28925]=61;
cos[28926]=61;
cos[28927]=61;
cos[28928]=61;
cos[28929]=61;
cos[28930]=61;
cos[28931]=61;
cos[28932]=61;
cos[28933]=61;
cos[28934]=61;
cos[28935]=61;
cos[28936]=61;
cos[28937]=61;
cos[28938]=61;
cos[28939]=61;
cos[28940]=61;
cos[28941]=61;
cos[28942]=61;
cos[28943]=62;
cos[28944]=62;
cos[28945]=62;
cos[28946]=62;
cos[28947]=62;
cos[28948]=62;
cos[28949]=62;
cos[28950]=62;
cos[28951]=62;
cos[28952]=62;
cos[28953]=62;
cos[28954]=62;
cos[28955]=62;
cos[28956]=62;
cos[28957]=62;
cos[28958]=62;
cos[28959]=62;
cos[28960]=62;
cos[28961]=62;
cos[28962]=62;
cos[28963]=62;
cos[28964]=62;
cos[28965]=62;
cos[28966]=62;
cos[28967]=62;
cos[28968]=62;
cos[28969]=62;
cos[28970]=62;
cos[28971]=62;
cos[28972]=62;
cos[28973]=62;
cos[28974]=62;
cos[28975]=62;
cos[28976]=63;
cos[28977]=63;
cos[28978]=63;
cos[28979]=63;
cos[28980]=63;
cos[28981]=63;
cos[28982]=63;
cos[28983]=63;
cos[28984]=63;
cos[28985]=63;
cos[28986]=63;
cos[28987]=63;
cos[28988]=63;
cos[28989]=63;
cos[28990]=63;
cos[28991]=63;
cos[28992]=63;
cos[28993]=63;
cos[28994]=63;
cos[28995]=63;
cos[28996]=63;
cos[28997]=63;
cos[28998]=63;
cos[28999]=63;
cos[29000]=63;
cos[29001]=63;
cos[29002]=63;
cos[29003]=63;
cos[29004]=63;
cos[29005]=63;
cos[29006]=63;
cos[29007]=63;
cos[29008]=63;
cos[29009]=63;
cos[29010]=63;
cos[29011]=64;
cos[29012]=64;
cos[29013]=64;
cos[29014]=64;
cos[29015]=64;
cos[29016]=64;
cos[29017]=64;
cos[29018]=64;
cos[29019]=64;
cos[29020]=64;
cos[29021]=64;
cos[29022]=64;
cos[29023]=64;
cos[29024]=64;
cos[29025]=64;
cos[29026]=64;
cos[29027]=64;
cos[29028]=64;
cos[29029]=64;
cos[29030]=64;
cos[29031]=64;
cos[29032]=64;
cos[29033]=64;
cos[29034]=64;
cos[29035]=64;
cos[29036]=64;
cos[29037]=64;
cos[29038]=64;
cos[29039]=64;
cos[29040]=64;
cos[29041]=64;
cos[29042]=64;
cos[29043]=64;
cos[29044]=64;
cos[29045]=64;
cos[29046]=65;
cos[29047]=65;
cos[29048]=65;
cos[29049]=65;
cos[29050]=65;
cos[29051]=65;
cos[29052]=65;
cos[29053]=65;
cos[29054]=65;
cos[29055]=65;
cos[29056]=65;
cos[29057]=65;
cos[29058]=65;
cos[29059]=65;
cos[29060]=65;
cos[29061]=65;
cos[29062]=65;
cos[29063]=65;
cos[29064]=65;
cos[29065]=65;
cos[29066]=65;
cos[29067]=65;
cos[29068]=65;
cos[29069]=65;
cos[29070]=65;
cos[29071]=65;
cos[29072]=65;
cos[29073]=65;
cos[29074]=65;
cos[29075]=65;
cos[29076]=65;
cos[29077]=65;
cos[29078]=65;
cos[29079]=65;
cos[29080]=65;
cos[29081]=65;
cos[29082]=65;
cos[29083]=66;
cos[29084]=66;
cos[29085]=66;
cos[29086]=66;
cos[29087]=66;
cos[29088]=66;
cos[29089]=66;
cos[29090]=66;
cos[29091]=66;
cos[29092]=66;
cos[29093]=66;
cos[29094]=66;
cos[29095]=66;
cos[29096]=66;
cos[29097]=66;
cos[29098]=66;
cos[29099]=66;
cos[29100]=66;
cos[29101]=66;
cos[29102]=66;
cos[29103]=66;
cos[29104]=66;
cos[29105]=66;
cos[29106]=66;
cos[29107]=66;
cos[29108]=66;
cos[29109]=66;
cos[29110]=66;
cos[29111]=66;
cos[29112]=66;
cos[29113]=66;
cos[29114]=66;
cos[29115]=66;
cos[29116]=66;
cos[29117]=66;
cos[29118]=66;
cos[29119]=66;
cos[29120]=66;
cos[29121]=67;
cos[29122]=67;
cos[29123]=67;
cos[29124]=67;
cos[29125]=67;
cos[29126]=67;
cos[29127]=67;
cos[29128]=67;
cos[29129]=67;
cos[29130]=67;
cos[29131]=67;
cos[29132]=67;
cos[29133]=67;
cos[29134]=67;
cos[29135]=67;
cos[29136]=67;
cos[29137]=67;
cos[29138]=67;
cos[29139]=67;
cos[29140]=67;
cos[29141]=67;
cos[29142]=67;
cos[29143]=67;
cos[29144]=67;
cos[29145]=67;
cos[29146]=67;
cos[29147]=67;
cos[29148]=67;
cos[29149]=67;
cos[29150]=67;
cos[29151]=67;
cos[29152]=67;
cos[29153]=67;
cos[29154]=67;
cos[29155]=67;
cos[29156]=67;
cos[29157]=67;
cos[29158]=67;
cos[29159]=67;
cos[29160]=67;
cos[29161]=68;
cos[29162]=68;
cos[29163]=68;
cos[29164]=68;
cos[29165]=68;
cos[29166]=68;
cos[29167]=68;
cos[29168]=68;
cos[29169]=68;
cos[29170]=68;
cos[29171]=68;
cos[29172]=68;
cos[29173]=68;
cos[29174]=68;
cos[29175]=68;
cos[29176]=68;
cos[29177]=68;
cos[29178]=68;
cos[29179]=68;
cos[29180]=68;
cos[29181]=68;
cos[29182]=68;
cos[29183]=68;
cos[29184]=68;
cos[29185]=68;
cos[29186]=68;
cos[29187]=68;
cos[29188]=68;
cos[29189]=68;
cos[29190]=68;
cos[29191]=68;
cos[29192]=68;
cos[29193]=68;
cos[29194]=68;
cos[29195]=68;
cos[29196]=68;
cos[29197]=68;
cos[29198]=68;
cos[29199]=68;
cos[29200]=68;
cos[29201]=68;
cos[29202]=69;
cos[29203]=69;
cos[29204]=69;
cos[29205]=69;
cos[29206]=69;
cos[29207]=69;
cos[29208]=69;
cos[29209]=69;
cos[29210]=69;
cos[29211]=69;
cos[29212]=69;
cos[29213]=69;
cos[29214]=69;
cos[29215]=69;
cos[29216]=69;
cos[29217]=69;
cos[29218]=69;
cos[29219]=69;
cos[29220]=69;
cos[29221]=69;
cos[29222]=69;
cos[29223]=69;
cos[29224]=69;
cos[29225]=69;
cos[29226]=69;
cos[29227]=69;
cos[29228]=69;
cos[29229]=69;
cos[29230]=69;
cos[29231]=69;
cos[29232]=69;
cos[29233]=69;
cos[29234]=69;
cos[29235]=69;
cos[29236]=69;
cos[29237]=69;
cos[29238]=69;
cos[29239]=69;
cos[29240]=69;
cos[29241]=69;
cos[29242]=69;
cos[29243]=69;
cos[29244]=69;
cos[29245]=69;
cos[29246]=70;
cos[29247]=70;
cos[29248]=70;
cos[29249]=70;
cos[29250]=70;
cos[29251]=70;
cos[29252]=70;
cos[29253]=70;
cos[29254]=70;
cos[29255]=70;
cos[29256]=70;
cos[29257]=70;
cos[29258]=70;
cos[29259]=70;
cos[29260]=70;
cos[29261]=70;
cos[29262]=70;
cos[29263]=70;
cos[29264]=70;
cos[29265]=70;
cos[29266]=70;
cos[29267]=70;
cos[29268]=70;
cos[29269]=70;
cos[29270]=70;
cos[29271]=70;
cos[29272]=70;
cos[29273]=70;
cos[29274]=70;
cos[29275]=70;
cos[29276]=70;
cos[29277]=70;
cos[29278]=70;
cos[29279]=70;
cos[29280]=70;
cos[29281]=70;
cos[29282]=70;
cos[29283]=70;
cos[29284]=70;
cos[29285]=70;
cos[29286]=70;
cos[29287]=70;
cos[29288]=70;
cos[29289]=70;
cos[29290]=70;
cos[29291]=71;
cos[29292]=71;
cos[29293]=71;
cos[29294]=71;
cos[29295]=71;
cos[29296]=71;
cos[29297]=71;
cos[29298]=71;
cos[29299]=71;
cos[29300]=71;
cos[29301]=71;
cos[29302]=71;
cos[29303]=71;
cos[29304]=71;
cos[29305]=71;
cos[29306]=71;
cos[29307]=71;
cos[29308]=71;
cos[29309]=71;
cos[29310]=71;
cos[29311]=71;
cos[29312]=71;
cos[29313]=71;
cos[29314]=71;
cos[29315]=71;
cos[29316]=71;
cos[29317]=71;
cos[29318]=71;
cos[29319]=71;
cos[29320]=71;
cos[29321]=71;
cos[29322]=71;
cos[29323]=71;
cos[29324]=71;
cos[29325]=71;
cos[29326]=71;
cos[29327]=71;
cos[29328]=71;
cos[29329]=71;
cos[29330]=71;
cos[29331]=71;
cos[29332]=71;
cos[29333]=71;
cos[29334]=71;
cos[29335]=71;
cos[29336]=71;
cos[29337]=71;
cos[29338]=71;
cos[29339]=71;
cos[29340]=72;
cos[29341]=72;
cos[29342]=72;
cos[29343]=72;
cos[29344]=72;
cos[29345]=72;
cos[29346]=72;
cos[29347]=72;
cos[29348]=72;
cos[29349]=72;
cos[29350]=72;
cos[29351]=72;
cos[29352]=72;
cos[29353]=72;
cos[29354]=72;
cos[29355]=72;
cos[29356]=72;
cos[29357]=72;
cos[29358]=72;
cos[29359]=72;
cos[29360]=72;
cos[29361]=72;
cos[29362]=72;
cos[29363]=72;
cos[29364]=72;
cos[29365]=72;
cos[29366]=72;
cos[29367]=72;
cos[29368]=72;
cos[29369]=72;
cos[29370]=72;
cos[29371]=72;
cos[29372]=72;
cos[29373]=72;
cos[29374]=72;
cos[29375]=72;
cos[29376]=72;
cos[29377]=72;
cos[29378]=72;
cos[29379]=72;
cos[29380]=72;
cos[29381]=72;
cos[29382]=72;
cos[29383]=72;
cos[29384]=72;
cos[29385]=72;
cos[29386]=72;
cos[29387]=72;
cos[29388]=72;
cos[29389]=72;
cos[29390]=72;
cos[29391]=72;
cos[29392]=72;
cos[29393]=73;
cos[29394]=73;
cos[29395]=73;
cos[29396]=73;
cos[29397]=73;
cos[29398]=73;
cos[29399]=73;
cos[29400]=73;
cos[29401]=73;
cos[29402]=73;
cos[29403]=73;
cos[29404]=73;
cos[29405]=73;
cos[29406]=73;
cos[29407]=73;
cos[29408]=73;
cos[29409]=73;
cos[29410]=73;
cos[29411]=73;
cos[29412]=73;
cos[29413]=73;
cos[29414]=73;
cos[29415]=73;
cos[29416]=73;
cos[29417]=73;
cos[29418]=73;
cos[29419]=73;
cos[29420]=73;
cos[29421]=73;
cos[29422]=73;
cos[29423]=73;
cos[29424]=73;
cos[29425]=73;
cos[29426]=73;
cos[29427]=73;
cos[29428]=73;
cos[29429]=73;
cos[29430]=73;
cos[29431]=73;
cos[29432]=73;
cos[29433]=73;
cos[29434]=73;
cos[29435]=73;
cos[29436]=73;
cos[29437]=73;
cos[29438]=73;
cos[29439]=73;
cos[29440]=73;
cos[29441]=73;
cos[29442]=73;
cos[29443]=73;
cos[29444]=73;
cos[29445]=73;
cos[29446]=73;
cos[29447]=73;
cos[29448]=73;
cos[29449]=73;
cos[29450]=74;
cos[29451]=74;
cos[29452]=74;
cos[29453]=74;
cos[29454]=74;
cos[29455]=74;
cos[29456]=74;
cos[29457]=74;
cos[29458]=74;
cos[29459]=74;
cos[29460]=74;
cos[29461]=74;
cos[29462]=74;
cos[29463]=74;
cos[29464]=74;
cos[29465]=74;
cos[29466]=74;
cos[29467]=74;
cos[29468]=74;
cos[29469]=74;
cos[29470]=74;
cos[29471]=74;
cos[29472]=74;
cos[29473]=74;
cos[29474]=74;
cos[29475]=74;
cos[29476]=74;
cos[29477]=74;
cos[29478]=74;
cos[29479]=74;
cos[29480]=74;
cos[29481]=74;
cos[29482]=74;
cos[29483]=74;
cos[29484]=74;
cos[29485]=74;
cos[29486]=74;
cos[29487]=74;
cos[29488]=74;
cos[29489]=74;
cos[29490]=74;
cos[29491]=74;
cos[29492]=74;
cos[29493]=74;
cos[29494]=74;
cos[29495]=74;
cos[29496]=74;
cos[29497]=74;
cos[29498]=74;
cos[29499]=74;
cos[29500]=74;
cos[29501]=74;
cos[29502]=74;
cos[29503]=74;
cos[29504]=74;
cos[29505]=74;
cos[29506]=74;
cos[29507]=74;
cos[29508]=74;
cos[29509]=74;
cos[29510]=74;
cos[29511]=74;
cos[29512]=74;
cos[29513]=74;
cos[29514]=75;
cos[29515]=75;
cos[29516]=75;
cos[29517]=75;
cos[29518]=75;
cos[29519]=75;
cos[29520]=75;
cos[29521]=75;
cos[29522]=75;
cos[29523]=75;
cos[29524]=75;
cos[29525]=75;
cos[29526]=75;
cos[29527]=75;
cos[29528]=75;
cos[29529]=75;
cos[29530]=75;
cos[29531]=75;
cos[29532]=75;
cos[29533]=75;
cos[29534]=75;
cos[29535]=75;
cos[29536]=75;
cos[29537]=75;
cos[29538]=75;
cos[29539]=75;
cos[29540]=75;
cos[29541]=75;
cos[29542]=75;
cos[29543]=75;
cos[29544]=75;
cos[29545]=75;
cos[29546]=75;
cos[29547]=75;
cos[29548]=75;
cos[29549]=75;
cos[29550]=75;
cos[29551]=75;
cos[29552]=75;
cos[29553]=75;
cos[29554]=75;
cos[29555]=75;
cos[29556]=75;
cos[29557]=75;
cos[29558]=75;
cos[29559]=75;
cos[29560]=75;
cos[29561]=75;
cos[29562]=75;
cos[29563]=75;
cos[29564]=75;
cos[29565]=75;
cos[29566]=75;
cos[29567]=75;
cos[29568]=75;
cos[29569]=75;
cos[29570]=75;
cos[29571]=75;
cos[29572]=75;
cos[29573]=75;
cos[29574]=75;
cos[29575]=75;
cos[29576]=75;
cos[29577]=75;
cos[29578]=75;
cos[29579]=75;
cos[29580]=75;
cos[29581]=75;
cos[29582]=75;
cos[29583]=75;
cos[29584]=75;
cos[29585]=75;
cos[29586]=75;
cos[29587]=76;
cos[29588]=76;
cos[29589]=76;
cos[29590]=76;
cos[29591]=76;
cos[29592]=76;
cos[29593]=76;
cos[29594]=76;
cos[29595]=76;
cos[29596]=76;
cos[29597]=76;
cos[29598]=76;
cos[29599]=76;
cos[29600]=76;
cos[29601]=76;
cos[29602]=76;
cos[29603]=76;
cos[29604]=76;
cos[29605]=76;
cos[29606]=76;
cos[29607]=76;
cos[29608]=76;
cos[29609]=76;
cos[29610]=76;
cos[29611]=76;
cos[29612]=76;
cos[29613]=76;
cos[29614]=76;
cos[29615]=76;
cos[29616]=76;
cos[29617]=76;
cos[29618]=76;
cos[29619]=76;
cos[29620]=76;
cos[29621]=76;
cos[29622]=76;
cos[29623]=76;
cos[29624]=76;
cos[29625]=76;
cos[29626]=76;
cos[29627]=76;
cos[29628]=76;
cos[29629]=76;
cos[29630]=76;
cos[29631]=76;
cos[29632]=76;
cos[29633]=76;
cos[29634]=76;
cos[29635]=76;
cos[29636]=76;
cos[29637]=76;
cos[29638]=76;
cos[29639]=76;
cos[29640]=76;
cos[29641]=76;
cos[29642]=76;
cos[29643]=76;
cos[29644]=76;
cos[29645]=76;
cos[29646]=76;
cos[29647]=76;
cos[29648]=76;
cos[29649]=76;
cos[29650]=76;
cos[29651]=76;
cos[29652]=76;
cos[29653]=76;
cos[29654]=76;
cos[29655]=76;
cos[29656]=76;
cos[29657]=76;
cos[29658]=76;
cos[29659]=76;
cos[29660]=76;
cos[29661]=76;
cos[29662]=76;
cos[29663]=76;
cos[29664]=76;
cos[29665]=76;
cos[29666]=76;
cos[29667]=76;
cos[29668]=76;
cos[29669]=76;
cos[29670]=76;
cos[29671]=76;
cos[29672]=76;
cos[29673]=76;
cos[29674]=76;
cos[29675]=77;
cos[29676]=77;
cos[29677]=77;
cos[29678]=77;
cos[29679]=77;
cos[29680]=77;
cos[29681]=77;
cos[29682]=77;
cos[29683]=77;
cos[29684]=77;
cos[29685]=77;
cos[29686]=77;
cos[29687]=77;
cos[29688]=77;
cos[29689]=77;
cos[29690]=77;
cos[29691]=77;
cos[29692]=77;
cos[29693]=77;
cos[29694]=77;
cos[29695]=77;
cos[29696]=77;
cos[29697]=77;
cos[29698]=77;
cos[29699]=77;
cos[29700]=77;
cos[29701]=77;
cos[29702]=77;
cos[29703]=77;
cos[29704]=77;
cos[29705]=77;
cos[29706]=77;
cos[29707]=77;
cos[29708]=77;
cos[29709]=77;
cos[29710]=77;
cos[29711]=77;
cos[29712]=77;
cos[29713]=77;
cos[29714]=77;
cos[29715]=77;
cos[29716]=77;
cos[29717]=77;
cos[29718]=77;
cos[29719]=77;
cos[29720]=77;
cos[29721]=77;
cos[29722]=77;
cos[29723]=77;
cos[29724]=77;
cos[29725]=77;
cos[29726]=77;
cos[29727]=77;
cos[29728]=77;
cos[29729]=77;
cos[29730]=77;
cos[29731]=77;
cos[29732]=77;
cos[29733]=77;
cos[29734]=77;
cos[29735]=77;
cos[29736]=77;
cos[29737]=77;
cos[29738]=77;
cos[29739]=77;
cos[29740]=77;
cos[29741]=77;
cos[29742]=77;
cos[29743]=77;
cos[29744]=77;
cos[29745]=77;
cos[29746]=77;
cos[29747]=77;
cos[29748]=77;
cos[29749]=77;
cos[29750]=77;
cos[29751]=77;
cos[29752]=77;
cos[29753]=77;
cos[29754]=77;
cos[29755]=77;
cos[29756]=77;
cos[29757]=77;
cos[29758]=77;
cos[29759]=77;
cos[29760]=77;
cos[29761]=77;
cos[29762]=77;
cos[29763]=77;
cos[29764]=77;
cos[29765]=77;
cos[29766]=77;
cos[29767]=77;
cos[29768]=77;
cos[29769]=77;
cos[29770]=77;
cos[29771]=77;
cos[29772]=77;
cos[29773]=77;
cos[29774]=77;
cos[29775]=77;
cos[29776]=77;
cos[29777]=77;
cos[29778]=77;
cos[29779]=77;
cos[29780]=77;
cos[29781]=77;
cos[29782]=77;
cos[29783]=77;
cos[29784]=77;
cos[29785]=77;
cos[29786]=77;
cos[29787]=77;
cos[29788]=77;
cos[29789]=77;
cos[29790]=77;
cos[29791]=77;
cos[29792]=77;
cos[29793]=77;
cos[29794]=77;
cos[29795]=77;
cos[29796]=77;
cos[29797]=77;
cos[29798]=77;
cos[29799]=78;
cos[29800]=78;
cos[29801]=78;
cos[29802]=78;
cos[29803]=78;
cos[29804]=78;
cos[29805]=78;
cos[29806]=78;
cos[29807]=78;
cos[29808]=78;
cos[29809]=78;
cos[29810]=78;
cos[29811]=78;
cos[29812]=78;
cos[29813]=78;
cos[29814]=78;
cos[29815]=78;
cos[29816]=78;
cos[29817]=78;
cos[29818]=78;
cos[29819]=78;
cos[29820]=78;
cos[29821]=78;
cos[29822]=78;
cos[29823]=78;
cos[29824]=78;
cos[29825]=78;
cos[29826]=78;
cos[29827]=78;
cos[29828]=78;
cos[29829]=78;
cos[29830]=78;
cos[29831]=78;
cos[29832]=78;
cos[29833]=78;
cos[29834]=78;
cos[29835]=78;
cos[29836]=78;
cos[29837]=78;
cos[29838]=78;
cos[29839]=78;
cos[29840]=78;
cos[29841]=78;
cos[29842]=78;
cos[29843]=78;
cos[29844]=78;
cos[29845]=78;
cos[29846]=78;
cos[29847]=78;
cos[29848]=78;
cos[29849]=78;
cos[29850]=78;
cos[29851]=78;
cos[29852]=78;
cos[29853]=78;
cos[29854]=78;
cos[29855]=78;
cos[29856]=78;
cos[29857]=78;
cos[29858]=78;
cos[29859]=78;
cos[29860]=78;
cos[29861]=78;
cos[29862]=78;
cos[29863]=78;
cos[29864]=78;
cos[29865]=78;
cos[29866]=78;
cos[29867]=78;
cos[29868]=78;
cos[29869]=78;
cos[29870]=78;
cos[29871]=78;
cos[29872]=78;
cos[29873]=78;
cos[29874]=78;
cos[29875]=78;
cos[29876]=78;
cos[29877]=78;
cos[29878]=78;
cos[29879]=78;
cos[29880]=78;
cos[29881]=78;
cos[29882]=78;
cos[29883]=78;
cos[29884]=78;
cos[29885]=78;
cos[29886]=78;
cos[29887]=78;
cos[29888]=78;
cos[29889]=78;
cos[29890]=78;
cos[29891]=78;
cos[29892]=78;
cos[29893]=78;
cos[29894]=78;
cos[29895]=78;
cos[29896]=78;
cos[29897]=78;
cos[29898]=78;
cos[29899]=78;
cos[29900]=78;
cos[29901]=78;
cos[29902]=78;
cos[29903]=78;
cos[29904]=78;
cos[29905]=78;
cos[29906]=78;
cos[29907]=78;
cos[29908]=78;
cos[29909]=78;
cos[29910]=78;
cos[29911]=78;
cos[29912]=78;
cos[29913]=78;
cos[29914]=78;
cos[29915]=78;
cos[29916]=78;
cos[29917]=78;
cos[29918]=78;
cos[29919]=78;
cos[29920]=78;
cos[29921]=78;
cos[29922]=78;
cos[29923]=78;
cos[29924]=78;
cos[29925]=78;
cos[29926]=78;
cos[29927]=78;
cos[29928]=78;
cos[29929]=78;
cos[29930]=78;
cos[29931]=78;
cos[29932]=78;
cos[29933]=78;
cos[29934]=78;
cos[29935]=78;
cos[29936]=78;
cos[29937]=78;
cos[29938]=78;
cos[29939]=78;
cos[29940]=78;
cos[29941]=78;
cos[29942]=78;
cos[29943]=78;
cos[29944]=78;
cos[29945]=78;
cos[29946]=78;
cos[29947]=78;
cos[29948]=78;
cos[29949]=78;
cos[29950]=78;
cos[29951]=78;
cos[29952]=78;
cos[29953]=78;
cos[29954]=78;
cos[29955]=78;
cos[29956]=78;
cos[29957]=78;
cos[29958]=78;
cos[29959]=78;
cos[29960]=78;
cos[29961]=78;
cos[29962]=78;
cos[29963]=78;
cos[29964]=78;
cos[29965]=78;
cos[29966]=78;
cos[29967]=78;
cos[29968]=78;
cos[29969]=78;
cos[29970]=78;
cos[29971]=78;
cos[29972]=78;
cos[29973]=78;
cos[29974]=78;
cos[29975]=78;
cos[29976]=78;
cos[29977]=78;
cos[29978]=78;
cos[29979]=78;
cos[29980]=78;
cos[29981]=78;
cos[29982]=78;
cos[29983]=78;
cos[29984]=78;
cos[29985]=78;
cos[29986]=78;
cos[29987]=78;
cos[29988]=78;
cos[29989]=78;
cos[29990]=78;
cos[29991]=78;
cos[29992]=78;
cos[29993]=78;
cos[29994]=78;
cos[29995]=78;
cos[29996]=78;
cos[29997]=78;
cos[29998]=78;
cos[29999]=78;
cos[30000]=78;
cos[30001]=78;
cos[30002]=78;
cos[30003]=78;
cos[30004]=78;
cos[30005]=78;
cos[30006]=78;
cos[30007]=78;
cos[30008]=78;
cos[30009]=78;
cos[30010]=78;
cos[30011]=78;
cos[30012]=78;
cos[30013]=78;
cos[30014]=78;
cos[30015]=78;
cos[30016]=78;
cos[30017]=78;
cos[30018]=78;
cos[30019]=78;
cos[30020]=78;
cos[30021]=78;
cos[30022]=78;
cos[30023]=78;
cos[30024]=78;
cos[30025]=78;
cos[30026]=78;
cos[30027]=78;
cos[30028]=78;
cos[30029]=78;
cos[30030]=78;
cos[30031]=78;
cos[30032]=78;
cos[30033]=78;
cos[30034]=78;
cos[30035]=78;
cos[30036]=78;
cos[30037]=78;
cos[30038]=78;
cos[30039]=78;
cos[30040]=78;
cos[30041]=78;
cos[30042]=78;
cos[30043]=78;
cos[30044]=78;
cos[30045]=78;
cos[30046]=78;
cos[30047]=78;
cos[30048]=78;
cos[30049]=78;
cos[30050]=78;
cos[30051]=78;
cos[30052]=78;
cos[30053]=78;
cos[30054]=78;
cos[30055]=78;
cos[30056]=78;
cos[30057]=78;
cos[30058]=78;
cos[30059]=78;
cos[30060]=78;
cos[30061]=78;
cos[30062]=78;
cos[30063]=78;
cos[30064]=78;
cos[30065]=78;
cos[30066]=78;
cos[30067]=78;
cos[30068]=78;
cos[30069]=78;
cos[30070]=78;
cos[30071]=78;
cos[30072]=78;
cos[30073]=78;
cos[30074]=78;
cos[30075]=78;
cos[30076]=78;
cos[30077]=78;
cos[30078]=78;
cos[30079]=78;
cos[30080]=78;
cos[30081]=78;
cos[30082]=78;
cos[30083]=78;
cos[30084]=78;
cos[30085]=78;
cos[30086]=78;
cos[30087]=78;
cos[30088]=78;
cos[30089]=78;
cos[30090]=78;
cos[30091]=78;
cos[30092]=78;
cos[30093]=78;
cos[30094]=78;
cos[30095]=78;
cos[30096]=78;
cos[30097]=78;
cos[30098]=78;
cos[30099]=78;
cos[30100]=78;
cos[30101]=78;
cos[30102]=78;
cos[30103]=78;
cos[30104]=78;
cos[30105]=78;
cos[30106]=78;
cos[30107]=78;
cos[30108]=78;
cos[30109]=78;
cos[30110]=78;
cos[30111]=78;
cos[30112]=78;
cos[30113]=78;
cos[30114]=78;
cos[30115]=78;
cos[30116]=78;
cos[30117]=78;
cos[30118]=78;
cos[30119]=78;
cos[30120]=78;
cos[30121]=78;
cos[30122]=78;
cos[30123]=78;
cos[30124]=78;
cos[30125]=78;
cos[30126]=78;
cos[30127]=78;
cos[30128]=78;
cos[30129]=78;
cos[30130]=78;
cos[30131]=78;
cos[30132]=78;
cos[30133]=78;
cos[30134]=78;
cos[30135]=78;
cos[30136]=78;
cos[30137]=78;
cos[30138]=78;
cos[30139]=78;
cos[30140]=78;
cos[30141]=78;
cos[30142]=78;
cos[30143]=78;
cos[30144]=78;
cos[30145]=78;
cos[30146]=78;
cos[30147]=78;
cos[30148]=78;
cos[30149]=78;
cos[30150]=78;
cos[30151]=78;
cos[30152]=78;
cos[30153]=78;
cos[30154]=78;
cos[30155]=78;
cos[30156]=78;
cos[30157]=78;
cos[30158]=78;
cos[30159]=78;
cos[30160]=78;
cos[30161]=78;
cos[30162]=78;
cos[30163]=78;
cos[30164]=78;
cos[30165]=78;
cos[30166]=78;
cos[30167]=78;
cos[30168]=78;
cos[30169]=78;
cos[30170]=78;
cos[30171]=78;
cos[30172]=78;
cos[30173]=78;
cos[30174]=78;
cos[30175]=78;
cos[30176]=78;
cos[30177]=78;
cos[30178]=78;
cos[30179]=78;
cos[30180]=78;
cos[30181]=78;
cos[30182]=78;
cos[30183]=78;
cos[30184]=78;
cos[30185]=78;
cos[30186]=78;
cos[30187]=78;
cos[30188]=78;
cos[30189]=78;
cos[30190]=78;
cos[30191]=78;
cos[30192]=78;
cos[30193]=78;
cos[30194]=78;
cos[30195]=78;
cos[30196]=78;
cos[30197]=78;
cos[30198]=78;
cos[30199]=78;
cos[30200]=78;
cos[30201]=78;
cos[30202]=77;
cos[30203]=77;
cos[30204]=77;
cos[30205]=77;
cos[30206]=77;
cos[30207]=77;
cos[30208]=77;
cos[30209]=77;
cos[30210]=77;
cos[30211]=77;
cos[30212]=77;
cos[30213]=77;
cos[30214]=77;
cos[30215]=77;
cos[30216]=77;
cos[30217]=77;
cos[30218]=77;
cos[30219]=77;
cos[30220]=77;
cos[30221]=77;
cos[30222]=77;
cos[30223]=77;
cos[30224]=77;
cos[30225]=77;
cos[30226]=77;
cos[30227]=77;
cos[30228]=77;
cos[30229]=77;
cos[30230]=77;
cos[30231]=77;
cos[30232]=77;
cos[30233]=77;
cos[30234]=77;
cos[30235]=77;
cos[30236]=77;
cos[30237]=77;
cos[30238]=77;
cos[30239]=77;
cos[30240]=77;
cos[30241]=77;
cos[30242]=77;
cos[30243]=77;
cos[30244]=77;
cos[30245]=77;
cos[30246]=77;
cos[30247]=77;
cos[30248]=77;
cos[30249]=77;
cos[30250]=77;
cos[30251]=77;
cos[30252]=77;
cos[30253]=77;
cos[30254]=77;
cos[30255]=77;
cos[30256]=77;
cos[30257]=77;
cos[30258]=77;
cos[30259]=77;
cos[30260]=77;
cos[30261]=77;
cos[30262]=77;
cos[30263]=77;
cos[30264]=77;
cos[30265]=77;
cos[30266]=77;
cos[30267]=77;
cos[30268]=77;
cos[30269]=77;
cos[30270]=77;
cos[30271]=77;
cos[30272]=77;
cos[30273]=77;
cos[30274]=77;
cos[30275]=77;
cos[30276]=77;
cos[30277]=77;
cos[30278]=77;
cos[30279]=77;
cos[30280]=77;
cos[30281]=77;
cos[30282]=77;
cos[30283]=77;
cos[30284]=77;
cos[30285]=77;
cos[30286]=77;
cos[30287]=77;
cos[30288]=77;
cos[30289]=77;
cos[30290]=77;
cos[30291]=77;
cos[30292]=77;
cos[30293]=77;
cos[30294]=77;
cos[30295]=77;
cos[30296]=77;
cos[30297]=77;
cos[30298]=77;
cos[30299]=77;
cos[30300]=77;
cos[30301]=77;
cos[30302]=77;
cos[30303]=77;
cos[30304]=77;
cos[30305]=77;
cos[30306]=77;
cos[30307]=77;
cos[30308]=77;
cos[30309]=77;
cos[30310]=77;
cos[30311]=77;
cos[30312]=77;
cos[30313]=77;
cos[30314]=77;
cos[30315]=77;
cos[30316]=77;
cos[30317]=77;
cos[30318]=77;
cos[30319]=77;
cos[30320]=77;
cos[30321]=77;
cos[30322]=77;
cos[30323]=77;
cos[30324]=77;
cos[30325]=77;
cos[30326]=76;
cos[30327]=76;
cos[30328]=76;
cos[30329]=76;
cos[30330]=76;
cos[30331]=76;
cos[30332]=76;
cos[30333]=76;
cos[30334]=76;
cos[30335]=76;
cos[30336]=76;
cos[30337]=76;
cos[30338]=76;
cos[30339]=76;
cos[30340]=76;
cos[30341]=76;
cos[30342]=76;
cos[30343]=76;
cos[30344]=76;
cos[30345]=76;
cos[30346]=76;
cos[30347]=76;
cos[30348]=76;
cos[30349]=76;
cos[30350]=76;
cos[30351]=76;
cos[30352]=76;
cos[30353]=76;
cos[30354]=76;
cos[30355]=76;
cos[30356]=76;
cos[30357]=76;
cos[30358]=76;
cos[30359]=76;
cos[30360]=76;
cos[30361]=76;
cos[30362]=76;
cos[30363]=76;
cos[30364]=76;
cos[30365]=76;
cos[30366]=76;
cos[30367]=76;
cos[30368]=76;
cos[30369]=76;
cos[30370]=76;
cos[30371]=76;
cos[30372]=76;
cos[30373]=76;
cos[30374]=76;
cos[30375]=76;
cos[30376]=76;
cos[30377]=76;
cos[30378]=76;
cos[30379]=76;
cos[30380]=76;
cos[30381]=76;
cos[30382]=76;
cos[30383]=76;
cos[30384]=76;
cos[30385]=76;
cos[30386]=76;
cos[30387]=76;
cos[30388]=76;
cos[30389]=76;
cos[30390]=76;
cos[30391]=76;
cos[30392]=76;
cos[30393]=76;
cos[30394]=76;
cos[30395]=76;
cos[30396]=76;
cos[30397]=76;
cos[30398]=76;
cos[30399]=76;
cos[30400]=76;
cos[30401]=76;
cos[30402]=76;
cos[30403]=76;
cos[30404]=76;
cos[30405]=76;
cos[30406]=76;
cos[30407]=76;
cos[30408]=76;
cos[30409]=76;
cos[30410]=76;
cos[30411]=76;
cos[30412]=76;
cos[30413]=76;
cos[30414]=75;
cos[30415]=75;
cos[30416]=75;
cos[30417]=75;
cos[30418]=75;
cos[30419]=75;
cos[30420]=75;
cos[30421]=75;
cos[30422]=75;
cos[30423]=75;
cos[30424]=75;
cos[30425]=75;
cos[30426]=75;
cos[30427]=75;
cos[30428]=75;
cos[30429]=75;
cos[30430]=75;
cos[30431]=75;
cos[30432]=75;
cos[30433]=75;
cos[30434]=75;
cos[30435]=75;
cos[30436]=75;
cos[30437]=75;
cos[30438]=75;
cos[30439]=75;
cos[30440]=75;
cos[30441]=75;
cos[30442]=75;
cos[30443]=75;
cos[30444]=75;
cos[30445]=75;
cos[30446]=75;
cos[30447]=75;
cos[30448]=75;
cos[30449]=75;
cos[30450]=75;
cos[30451]=75;
cos[30452]=75;
cos[30453]=75;
cos[30454]=75;
cos[30455]=75;
cos[30456]=75;
cos[30457]=75;
cos[30458]=75;
cos[30459]=75;
cos[30460]=75;
cos[30461]=75;
cos[30462]=75;
cos[30463]=75;
cos[30464]=75;
cos[30465]=75;
cos[30466]=75;
cos[30467]=75;
cos[30468]=75;
cos[30469]=75;
cos[30470]=75;
cos[30471]=75;
cos[30472]=75;
cos[30473]=75;
cos[30474]=75;
cos[30475]=75;
cos[30476]=75;
cos[30477]=75;
cos[30478]=75;
cos[30479]=75;
cos[30480]=75;
cos[30481]=75;
cos[30482]=75;
cos[30483]=75;
cos[30484]=75;
cos[30485]=75;
cos[30486]=75;
cos[30487]=74;
cos[30488]=74;
cos[30489]=74;
cos[30490]=74;
cos[30491]=74;
cos[30492]=74;
cos[30493]=74;
cos[30494]=74;
cos[30495]=74;
cos[30496]=74;
cos[30497]=74;
cos[30498]=74;
cos[30499]=74;
cos[30500]=74;
cos[30501]=74;
cos[30502]=74;
cos[30503]=74;
cos[30504]=74;
cos[30505]=74;
cos[30506]=74;
cos[30507]=74;
cos[30508]=74;
cos[30509]=74;
cos[30510]=74;
cos[30511]=74;
cos[30512]=74;
cos[30513]=74;
cos[30514]=74;
cos[30515]=74;
cos[30516]=74;
cos[30517]=74;
cos[30518]=74;
cos[30519]=74;
cos[30520]=74;
cos[30521]=74;
cos[30522]=74;
cos[30523]=74;
cos[30524]=74;
cos[30525]=74;
cos[30526]=74;
cos[30527]=74;
cos[30528]=74;
cos[30529]=74;
cos[30530]=74;
cos[30531]=74;
cos[30532]=74;
cos[30533]=74;
cos[30534]=74;
cos[30535]=74;
cos[30536]=74;
cos[30537]=74;
cos[30538]=74;
cos[30539]=74;
cos[30540]=74;
cos[30541]=74;
cos[30542]=74;
cos[30543]=74;
cos[30544]=74;
cos[30545]=74;
cos[30546]=74;
cos[30547]=74;
cos[30548]=74;
cos[30549]=74;
cos[30550]=74;
cos[30551]=73;
cos[30552]=73;
cos[30553]=73;
cos[30554]=73;
cos[30555]=73;
cos[30556]=73;
cos[30557]=73;
cos[30558]=73;
cos[30559]=73;
cos[30560]=73;
cos[30561]=73;
cos[30562]=73;
cos[30563]=73;
cos[30564]=73;
cos[30565]=73;
cos[30566]=73;
cos[30567]=73;
cos[30568]=73;
cos[30569]=73;
cos[30570]=73;
cos[30571]=73;
cos[30572]=73;
cos[30573]=73;
cos[30574]=73;
cos[30575]=73;
cos[30576]=73;
cos[30577]=73;
cos[30578]=73;
cos[30579]=73;
cos[30580]=73;
cos[30581]=73;
cos[30582]=73;
cos[30583]=73;
cos[30584]=73;
cos[30585]=73;
cos[30586]=73;
cos[30587]=73;
cos[30588]=73;
cos[30589]=73;
cos[30590]=73;
cos[30591]=73;
cos[30592]=73;
cos[30593]=73;
cos[30594]=73;
cos[30595]=73;
cos[30596]=73;
cos[30597]=73;
cos[30598]=73;
cos[30599]=73;
cos[30600]=73;
cos[30601]=73;
cos[30602]=73;
cos[30603]=73;
cos[30604]=73;
cos[30605]=73;
cos[30606]=73;
cos[30607]=73;
cos[30608]=72;
cos[30609]=72;
cos[30610]=72;
cos[30611]=72;
cos[30612]=72;
cos[30613]=72;
cos[30614]=72;
cos[30615]=72;
cos[30616]=72;
cos[30617]=72;
cos[30618]=72;
cos[30619]=72;
cos[30620]=72;
cos[30621]=72;
cos[30622]=72;
cos[30623]=72;
cos[30624]=72;
cos[30625]=72;
cos[30626]=72;
cos[30627]=72;
cos[30628]=72;
cos[30629]=72;
cos[30630]=72;
cos[30631]=72;
cos[30632]=72;
cos[30633]=72;
cos[30634]=72;
cos[30635]=72;
cos[30636]=72;
cos[30637]=72;
cos[30638]=72;
cos[30639]=72;
cos[30640]=72;
cos[30641]=72;
cos[30642]=72;
cos[30643]=72;
cos[30644]=72;
cos[30645]=72;
cos[30646]=72;
cos[30647]=72;
cos[30648]=72;
cos[30649]=72;
cos[30650]=72;
cos[30651]=72;
cos[30652]=72;
cos[30653]=72;
cos[30654]=72;
cos[30655]=72;
cos[30656]=72;
cos[30657]=72;
cos[30658]=72;
cos[30659]=72;
cos[30660]=72;
cos[30661]=71;
cos[30662]=71;
cos[30663]=71;
cos[30664]=71;
cos[30665]=71;
cos[30666]=71;
cos[30667]=71;
cos[30668]=71;
cos[30669]=71;
cos[30670]=71;
cos[30671]=71;
cos[30672]=71;
cos[30673]=71;
cos[30674]=71;
cos[30675]=71;
cos[30676]=71;
cos[30677]=71;
cos[30678]=71;
cos[30679]=71;
cos[30680]=71;
cos[30681]=71;
cos[30682]=71;
cos[30683]=71;
cos[30684]=71;
cos[30685]=71;
cos[30686]=71;
cos[30687]=71;
cos[30688]=71;
cos[30689]=71;
cos[30690]=71;
cos[30691]=71;
cos[30692]=71;
cos[30693]=71;
cos[30694]=71;
cos[30695]=71;
cos[30696]=71;
cos[30697]=71;
cos[30698]=71;
cos[30699]=71;
cos[30700]=71;
cos[30701]=71;
cos[30702]=71;
cos[30703]=71;
cos[30704]=71;
cos[30705]=71;
cos[30706]=71;
cos[30707]=71;
cos[30708]=71;
cos[30709]=71;
cos[30710]=70;
cos[30711]=70;
cos[30712]=70;
cos[30713]=70;
cos[30714]=70;
cos[30715]=70;
cos[30716]=70;
cos[30717]=70;
cos[30718]=70;
cos[30719]=70;
cos[30720]=70;
cos[30721]=70;
cos[30722]=70;
cos[30723]=70;
cos[30724]=70;
cos[30725]=70;
cos[30726]=70;
cos[30727]=70;
cos[30728]=70;
cos[30729]=70;
cos[30730]=70;
cos[30731]=70;
cos[30732]=70;
cos[30733]=70;
cos[30734]=70;
cos[30735]=70;
cos[30736]=70;
cos[30737]=70;
cos[30738]=70;
cos[30739]=70;
cos[30740]=70;
cos[30741]=70;
cos[30742]=70;
cos[30743]=70;
cos[30744]=70;
cos[30745]=70;
cos[30746]=70;
cos[30747]=70;
cos[30748]=70;
cos[30749]=70;
cos[30750]=70;
cos[30751]=70;
cos[30752]=70;
cos[30753]=70;
cos[30754]=70;
cos[30755]=69;
cos[30756]=69;
cos[30757]=69;
cos[30758]=69;
cos[30759]=69;
cos[30760]=69;
cos[30761]=69;
cos[30762]=69;
cos[30763]=69;
cos[30764]=69;
cos[30765]=69;
cos[30766]=69;
cos[30767]=69;
cos[30768]=69;
cos[30769]=69;
cos[30770]=69;
cos[30771]=69;
cos[30772]=69;
cos[30773]=69;
cos[30774]=69;
cos[30775]=69;
cos[30776]=69;
cos[30777]=69;
cos[30778]=69;
cos[30779]=69;
cos[30780]=69;
cos[30781]=69;
cos[30782]=69;
cos[30783]=69;
cos[30784]=69;
cos[30785]=69;
cos[30786]=69;
cos[30787]=69;
cos[30788]=69;
cos[30789]=69;
cos[30790]=69;
cos[30791]=69;
cos[30792]=69;
cos[30793]=69;
cos[30794]=69;
cos[30795]=69;
cos[30796]=69;
cos[30797]=69;
cos[30798]=69;
cos[30799]=68;
cos[30800]=68;
cos[30801]=68;
cos[30802]=68;
cos[30803]=68;
cos[30804]=68;
cos[30805]=68;
cos[30806]=68;
cos[30807]=68;
cos[30808]=68;
cos[30809]=68;
cos[30810]=68;
cos[30811]=68;
cos[30812]=68;
cos[30813]=68;
cos[30814]=68;
cos[30815]=68;
cos[30816]=68;
cos[30817]=68;
cos[30818]=68;
cos[30819]=68;
cos[30820]=68;
cos[30821]=68;
cos[30822]=68;
cos[30823]=68;
cos[30824]=68;
cos[30825]=68;
cos[30826]=68;
cos[30827]=68;
cos[30828]=68;
cos[30829]=68;
cos[30830]=68;
cos[30831]=68;
cos[30832]=68;
cos[30833]=68;
cos[30834]=68;
cos[30835]=68;
cos[30836]=68;
cos[30837]=68;
cos[30838]=68;
cos[30839]=68;
cos[30840]=67;
cos[30841]=67;
cos[30842]=67;
cos[30843]=67;
cos[30844]=67;
cos[30845]=67;
cos[30846]=67;
cos[30847]=67;
cos[30848]=67;
cos[30849]=67;
cos[30850]=67;
cos[30851]=67;
cos[30852]=67;
cos[30853]=67;
cos[30854]=67;
cos[30855]=67;
cos[30856]=67;
cos[30857]=67;
cos[30858]=67;
cos[30859]=67;
cos[30860]=67;
cos[30861]=67;
cos[30862]=67;
cos[30863]=67;
cos[30864]=67;
cos[30865]=67;
cos[30866]=67;
cos[30867]=67;
cos[30868]=67;
cos[30869]=67;
cos[30870]=67;
cos[30871]=67;
cos[30872]=67;
cos[30873]=67;
cos[30874]=67;
cos[30875]=67;
cos[30876]=67;
cos[30877]=67;
cos[30878]=67;
cos[30879]=67;
cos[30880]=66;
cos[30881]=66;
cos[30882]=66;
cos[30883]=66;
cos[30884]=66;
cos[30885]=66;
cos[30886]=66;
cos[30887]=66;
cos[30888]=66;
cos[30889]=66;
cos[30890]=66;
cos[30891]=66;
cos[30892]=66;
cos[30893]=66;
cos[30894]=66;
cos[30895]=66;
cos[30896]=66;
cos[30897]=66;
cos[30898]=66;
cos[30899]=66;
cos[30900]=66;
cos[30901]=66;
cos[30902]=66;
cos[30903]=66;
cos[30904]=66;
cos[30905]=66;
cos[30906]=66;
cos[30907]=66;
cos[30908]=66;
cos[30909]=66;
cos[30910]=66;
cos[30911]=66;
cos[30912]=66;
cos[30913]=66;
cos[30914]=66;
cos[30915]=66;
cos[30916]=66;
cos[30917]=66;
cos[30918]=65;
cos[30919]=65;
cos[30920]=65;
cos[30921]=65;
cos[30922]=65;
cos[30923]=65;
cos[30924]=65;
cos[30925]=65;
cos[30926]=65;
cos[30927]=65;
cos[30928]=65;
cos[30929]=65;
cos[30930]=65;
cos[30931]=65;
cos[30932]=65;
cos[30933]=65;
cos[30934]=65;
cos[30935]=65;
cos[30936]=65;
cos[30937]=65;
cos[30938]=65;
cos[30939]=65;
cos[30940]=65;
cos[30941]=65;
cos[30942]=65;
cos[30943]=65;
cos[30944]=65;
cos[30945]=65;
cos[30946]=65;
cos[30947]=65;
cos[30948]=65;
cos[30949]=65;
cos[30950]=65;
cos[30951]=65;
cos[30952]=65;
cos[30953]=65;
cos[30954]=65;
cos[30955]=64;
cos[30956]=64;
cos[30957]=64;
cos[30958]=64;
cos[30959]=64;
cos[30960]=64;
cos[30961]=64;
cos[30962]=64;
cos[30963]=64;
cos[30964]=64;
cos[30965]=64;
cos[30966]=64;
cos[30967]=64;
cos[30968]=64;
cos[30969]=64;
cos[30970]=64;
cos[30971]=64;
cos[30972]=64;
cos[30973]=64;
cos[30974]=64;
cos[30975]=64;
cos[30976]=64;
cos[30977]=64;
cos[30978]=64;
cos[30979]=64;
cos[30980]=64;
cos[30981]=64;
cos[30982]=64;
cos[30983]=64;
cos[30984]=64;
cos[30985]=64;
cos[30986]=64;
cos[30987]=64;
cos[30988]=64;
cos[30989]=64;
cos[30990]=63;
cos[30991]=63;
cos[30992]=63;
cos[30993]=63;
cos[30994]=63;
cos[30995]=63;
cos[30996]=63;
cos[30997]=63;
cos[30998]=63;
cos[30999]=63;
cos[31000]=63;
cos[31001]=63;
cos[31002]=63;
cos[31003]=63;
cos[31004]=63;
cos[31005]=63;
cos[31006]=63;
cos[31007]=63;
cos[31008]=63;
cos[31009]=63;
cos[31010]=63;
cos[31011]=63;
cos[31012]=63;
cos[31013]=63;
cos[31014]=63;
cos[31015]=63;
cos[31016]=63;
cos[31017]=63;
cos[31018]=63;
cos[31019]=63;
cos[31020]=63;
cos[31021]=63;
cos[31022]=63;
cos[31023]=63;
cos[31024]=63;
cos[31025]=62;
cos[31026]=62;
cos[31027]=62;
cos[31028]=62;
cos[31029]=62;
cos[31030]=62;
cos[31031]=62;
cos[31032]=62;
cos[31033]=62;
cos[31034]=62;
cos[31035]=62;
cos[31036]=62;
cos[31037]=62;
cos[31038]=62;
cos[31039]=62;
cos[31040]=62;
cos[31041]=62;
cos[31042]=62;
cos[31043]=62;
cos[31044]=62;
cos[31045]=62;
cos[31046]=62;
cos[31047]=62;
cos[31048]=62;
cos[31049]=62;
cos[31050]=62;
cos[31051]=62;
cos[31052]=62;
cos[31053]=62;
cos[31054]=62;
cos[31055]=62;
cos[31056]=62;
cos[31057]=62;
cos[31058]=61;
cos[31059]=61;
cos[31060]=61;
cos[31061]=61;
cos[31062]=61;
cos[31063]=61;
cos[31064]=61;
cos[31065]=61;
cos[31066]=61;
cos[31067]=61;
cos[31068]=61;
cos[31069]=61;
cos[31070]=61;
cos[31071]=61;
cos[31072]=61;
cos[31073]=61;
cos[31074]=61;
cos[31075]=61;
cos[31076]=61;
cos[31077]=61;
cos[31078]=61;
cos[31079]=61;
cos[31080]=61;
cos[31081]=61;
cos[31082]=61;
cos[31083]=61;
cos[31084]=61;
cos[31085]=61;
cos[31086]=61;
cos[31087]=61;
cos[31088]=61;
cos[31089]=61;
cos[31090]=61;
cos[31091]=60;
cos[31092]=60;
cos[31093]=60;
cos[31094]=60;
cos[31095]=60;
cos[31096]=60;
cos[31097]=60;
cos[31098]=60;
cos[31099]=60;
cos[31100]=60;
cos[31101]=60;
cos[31102]=60;
cos[31103]=60;
cos[31104]=60;
cos[31105]=60;
cos[31106]=60;
cos[31107]=60;
cos[31108]=60;
cos[31109]=60;
cos[31110]=60;
cos[31111]=60;
cos[31112]=60;
cos[31113]=60;
cos[31114]=60;
cos[31115]=60;
cos[31116]=60;
cos[31117]=60;
cos[31118]=60;
cos[31119]=60;
cos[31120]=60;
cos[31121]=60;
cos[31122]=60;
cos[31123]=59;
cos[31124]=59;
cos[31125]=59;
cos[31126]=59;
cos[31127]=59;
cos[31128]=59;
cos[31129]=59;
cos[31130]=59;
cos[31131]=59;
cos[31132]=59;
cos[31133]=59;
cos[31134]=59;
cos[31135]=59;
cos[31136]=59;
cos[31137]=59;
cos[31138]=59;
cos[31139]=59;
cos[31140]=59;
cos[31141]=59;
cos[31142]=59;
cos[31143]=59;
cos[31144]=59;
cos[31145]=59;
cos[31146]=59;
cos[31147]=59;
cos[31148]=59;
cos[31149]=59;
cos[31150]=59;
cos[31151]=59;
cos[31152]=59;
cos[31153]=59;
cos[31154]=58;
cos[31155]=58;
cos[31156]=58;
cos[31157]=58;
cos[31158]=58;
cos[31159]=58;
cos[31160]=58;
cos[31161]=58;
cos[31162]=58;
cos[31163]=58;
cos[31164]=58;
cos[31165]=58;
cos[31166]=58;
cos[31167]=58;
cos[31168]=58;
cos[31169]=58;
cos[31170]=58;
cos[31171]=58;
cos[31172]=58;
cos[31173]=58;
cos[31174]=58;
cos[31175]=58;
cos[31176]=58;
cos[31177]=58;
cos[31178]=58;
cos[31179]=58;
cos[31180]=58;
cos[31181]=58;
cos[31182]=58;
cos[31183]=58;
cos[31184]=57;
cos[31185]=57;
cos[31186]=57;
cos[31187]=57;
cos[31188]=57;
cos[31189]=57;
cos[31190]=57;
cos[31191]=57;
cos[31192]=57;
cos[31193]=57;
cos[31194]=57;
cos[31195]=57;
cos[31196]=57;
cos[31197]=57;
cos[31198]=57;
cos[31199]=57;
cos[31200]=57;
cos[31201]=57;
cos[31202]=57;
cos[31203]=57;
cos[31204]=57;
cos[31205]=57;
cos[31206]=57;
cos[31207]=57;
cos[31208]=57;
cos[31209]=57;
cos[31210]=57;
cos[31211]=57;
cos[31212]=57;
cos[31213]=57;
cos[31214]=56;
cos[31215]=56;
cos[31216]=56;
cos[31217]=56;
cos[31218]=56;
cos[31219]=56;
cos[31220]=56;
cos[31221]=56;
cos[31222]=56;
cos[31223]=56;
cos[31224]=56;
cos[31225]=56;
cos[31226]=56;
cos[31227]=56;
cos[31228]=56;
cos[31229]=56;
cos[31230]=56;
cos[31231]=56;
cos[31232]=56;
cos[31233]=56;
cos[31234]=56;
cos[31235]=56;
cos[31236]=56;
cos[31237]=56;
cos[31238]=56;
cos[31239]=56;
cos[31240]=56;
cos[31241]=56;
cos[31242]=56;
cos[31243]=55;
cos[31244]=55;
cos[31245]=55;
cos[31246]=55;
cos[31247]=55;
cos[31248]=55;
cos[31249]=55;
cos[31250]=55;
cos[31251]=55;
cos[31252]=55;
cos[31253]=55;
cos[31254]=55;
cos[31255]=55;
cos[31256]=55;
cos[31257]=55;
cos[31258]=55;
cos[31259]=55;
cos[31260]=55;
cos[31261]=55;
cos[31262]=55;
cos[31263]=55;
cos[31264]=55;
cos[31265]=55;
cos[31266]=55;
cos[31267]=55;
cos[31268]=55;
cos[31269]=55;
cos[31270]=55;
cos[31271]=55;
cos[31272]=54;
cos[31273]=54;
cos[31274]=54;
cos[31275]=54;
cos[31276]=54;
cos[31277]=54;
cos[31278]=54;
cos[31279]=54;
cos[31280]=54;
cos[31281]=54;
cos[31282]=54;
cos[31283]=54;
cos[31284]=54;
cos[31285]=54;
cos[31286]=54;
cos[31287]=54;
cos[31288]=54;
cos[31289]=54;
cos[31290]=54;
cos[31291]=54;
cos[31292]=54;
cos[31293]=54;
cos[31294]=54;
cos[31295]=54;
cos[31296]=54;
cos[31297]=54;
cos[31298]=54;
cos[31299]=54;
cos[31300]=53;
cos[31301]=53;
cos[31302]=53;
cos[31303]=53;
cos[31304]=53;
cos[31305]=53;
cos[31306]=53;
cos[31307]=53;
cos[31308]=53;
cos[31309]=53;
cos[31310]=53;
cos[31311]=53;
cos[31312]=53;
cos[31313]=53;
cos[31314]=53;
cos[31315]=53;
cos[31316]=53;
cos[31317]=53;
cos[31318]=53;
cos[31319]=53;
cos[31320]=53;
cos[31321]=53;
cos[31322]=53;
cos[31323]=53;
cos[31324]=53;
cos[31325]=53;
cos[31326]=53;
cos[31327]=53;
cos[31328]=52;
cos[31329]=52;
cos[31330]=52;
cos[31331]=52;
cos[31332]=52;
cos[31333]=52;
cos[31334]=52;
cos[31335]=52;
cos[31336]=52;
cos[31337]=52;
cos[31338]=52;
cos[31339]=52;
cos[31340]=52;
cos[31341]=52;
cos[31342]=52;
cos[31343]=52;
cos[31344]=52;
cos[31345]=52;
cos[31346]=52;
cos[31347]=52;
cos[31348]=52;
cos[31349]=52;
cos[31350]=52;
cos[31351]=52;
cos[31352]=52;
cos[31353]=52;
cos[31354]=52;
cos[31355]=51;
cos[31356]=51;
cos[31357]=51;
cos[31358]=51;
cos[31359]=51;
cos[31360]=51;
cos[31361]=51;
cos[31362]=51;
cos[31363]=51;
cos[31364]=51;
cos[31365]=51;
cos[31366]=51;
cos[31367]=51;
cos[31368]=51;
cos[31369]=51;
cos[31370]=51;
cos[31371]=51;
cos[31372]=51;
cos[31373]=51;
cos[31374]=51;
cos[31375]=51;
cos[31376]=51;
cos[31377]=51;
cos[31378]=51;
cos[31379]=51;
cos[31380]=51;
cos[31381]=51;
cos[31382]=50;
cos[31383]=50;
cos[31384]=50;
cos[31385]=50;
cos[31386]=50;
cos[31387]=50;
cos[31388]=50;
cos[31389]=50;
cos[31390]=50;
cos[31391]=50;
cos[31392]=50;
cos[31393]=50;
cos[31394]=50;
cos[31395]=50;
cos[31396]=50;
cos[31397]=50;
cos[31398]=50;
cos[31399]=50;
cos[31400]=50;
cos[31401]=50;
cos[31402]=50;
cos[31403]=50;
cos[31404]=50;
cos[31405]=50;
cos[31406]=50;
cos[31407]=50;
cos[31408]=49;
cos[31409]=49;
cos[31410]=49;
cos[31411]=49;
cos[31412]=49;
cos[31413]=49;
cos[31414]=49;
cos[31415]=49;
cos[31416]=49;
cos[31417]=49;
cos[31418]=49;
cos[31419]=49;
cos[31420]=49;
cos[31421]=49;
cos[31422]=49;
cos[31423]=49;
cos[31424]=49;
cos[31425]=49;
cos[31426]=49;
cos[31427]=49;
cos[31428]=49;
cos[31429]=49;
cos[31430]=49;
cos[31431]=49;
cos[31432]=49;
cos[31433]=49;
cos[31434]=49;
cos[31435]=48;
cos[31436]=48;
cos[31437]=48;
cos[31438]=48;
cos[31439]=48;
cos[31440]=48;
cos[31441]=48;
cos[31442]=48;
cos[31443]=48;
cos[31444]=48;
cos[31445]=48;
cos[31446]=48;
cos[31447]=48;
cos[31448]=48;
cos[31449]=48;
cos[31450]=48;
cos[31451]=48;
cos[31452]=48;
cos[31453]=48;
cos[31454]=48;
cos[31455]=48;
cos[31456]=48;
cos[31457]=48;
cos[31458]=48;
cos[31459]=48;
cos[31460]=47;
cos[31461]=47;
cos[31462]=47;
cos[31463]=47;
cos[31464]=47;
cos[31465]=47;
cos[31466]=47;
cos[31467]=47;
cos[31468]=47;
cos[31469]=47;
cos[31470]=47;
cos[31471]=47;
cos[31472]=47;
cos[31473]=47;
cos[31474]=47;
cos[31475]=47;
cos[31476]=47;
cos[31477]=47;
cos[31478]=47;
cos[31479]=47;
cos[31480]=47;
cos[31481]=47;
cos[31482]=47;
cos[31483]=47;
cos[31484]=47;
cos[31485]=47;
cos[31486]=46;
cos[31487]=46;
cos[31488]=46;
cos[31489]=46;
cos[31490]=46;
cos[31491]=46;
cos[31492]=46;
cos[31493]=46;
cos[31494]=46;
cos[31495]=46;
cos[31496]=46;
cos[31497]=46;
cos[31498]=46;
cos[31499]=46;
cos[31500]=46;
cos[31501]=46;
cos[31502]=46;
cos[31503]=46;
cos[31504]=46;
cos[31505]=46;
cos[31506]=46;
cos[31507]=46;
cos[31508]=46;
cos[31509]=46;
cos[31510]=46;
cos[31511]=45;
cos[31512]=45;
cos[31513]=45;
cos[31514]=45;
cos[31515]=45;
cos[31516]=45;
cos[31517]=45;
cos[31518]=45;
cos[31519]=45;
cos[31520]=45;
cos[31521]=45;
cos[31522]=45;
cos[31523]=45;
cos[31524]=45;
cos[31525]=45;
cos[31526]=45;
cos[31527]=45;
cos[31528]=45;
cos[31529]=45;
cos[31530]=45;
cos[31531]=45;
cos[31532]=45;
cos[31533]=45;
cos[31534]=45;
cos[31535]=45;
cos[31536]=44;
cos[31537]=44;
cos[31538]=44;
cos[31539]=44;
cos[31540]=44;
cos[31541]=44;
cos[31542]=44;
cos[31543]=44;
cos[31544]=44;
cos[31545]=44;
cos[31546]=44;
cos[31547]=44;
cos[31548]=44;
cos[31549]=44;
cos[31550]=44;
cos[31551]=44;
cos[31552]=44;
cos[31553]=44;
cos[31554]=44;
cos[31555]=44;
cos[31556]=44;
cos[31557]=44;
cos[31558]=44;
cos[31559]=44;
cos[31560]=44;
cos[31561]=43;
cos[31562]=43;
cos[31563]=43;
cos[31564]=43;
cos[31565]=43;
cos[31566]=43;
cos[31567]=43;
cos[31568]=43;
cos[31569]=43;
cos[31570]=43;
cos[31571]=43;
cos[31572]=43;
cos[31573]=43;
cos[31574]=43;
cos[31575]=43;
cos[31576]=43;
cos[31577]=43;
cos[31578]=43;
cos[31579]=43;
cos[31580]=43;
cos[31581]=43;
cos[31582]=43;
cos[31583]=43;
cos[31584]=43;
cos[31585]=42;
cos[31586]=42;
cos[31587]=42;
cos[31588]=42;
cos[31589]=42;
cos[31590]=42;
cos[31591]=42;
cos[31592]=42;
cos[31593]=42;
cos[31594]=42;
cos[31595]=42;
cos[31596]=42;
cos[31597]=42;
cos[31598]=42;
cos[31599]=42;
cos[31600]=42;
cos[31601]=42;
cos[31602]=42;
cos[31603]=42;
cos[31604]=42;
cos[31605]=42;
cos[31606]=42;
cos[31607]=42;
cos[31608]=42;
cos[31609]=41;
cos[31610]=41;
cos[31611]=41;
cos[31612]=41;
cos[31613]=41;
cos[31614]=41;
cos[31615]=41;
cos[31616]=41;
cos[31617]=41;
cos[31618]=41;
cos[31619]=41;
cos[31620]=41;
cos[31621]=41;
cos[31622]=41;
cos[31623]=41;
cos[31624]=41;
cos[31625]=41;
cos[31626]=41;
cos[31627]=41;
cos[31628]=41;
cos[31629]=41;
cos[31630]=41;
cos[31631]=41;
cos[31632]=41;
cos[31633]=40;
cos[31634]=40;
cos[31635]=40;
cos[31636]=40;
cos[31637]=40;
cos[31638]=40;
cos[31639]=40;
cos[31640]=40;
cos[31641]=40;
cos[31642]=40;
cos[31643]=40;
cos[31644]=40;
cos[31645]=40;
cos[31646]=40;
cos[31647]=40;
cos[31648]=40;
cos[31649]=40;
cos[31650]=40;
cos[31651]=40;
cos[31652]=40;
cos[31653]=40;
cos[31654]=40;
cos[31655]=40;
cos[31656]=40;
cos[31657]=39;
cos[31658]=39;
cos[31659]=39;
cos[31660]=39;
cos[31661]=39;
cos[31662]=39;
cos[31663]=39;
cos[31664]=39;
cos[31665]=39;
cos[31666]=39;
cos[31667]=39;
cos[31668]=39;
cos[31669]=39;
cos[31670]=39;
cos[31671]=39;
cos[31672]=39;
cos[31673]=39;
cos[31674]=39;
cos[31675]=39;
cos[31676]=39;
cos[31677]=39;
cos[31678]=39;
cos[31679]=39;
cos[31680]=38;
cos[31681]=38;
cos[31682]=38;
cos[31683]=38;
cos[31684]=38;
cos[31685]=38;
cos[31686]=38;
cos[31687]=38;
cos[31688]=38;
cos[31689]=38;
cos[31690]=38;
cos[31691]=38;
cos[31692]=38;
cos[31693]=38;
cos[31694]=38;
cos[31695]=38;
cos[31696]=38;
cos[31697]=38;
cos[31698]=38;
cos[31699]=38;
cos[31700]=38;
cos[31701]=38;
cos[31702]=38;
cos[31703]=38;
cos[31704]=37;
cos[31705]=37;
cos[31706]=37;
cos[31707]=37;
cos[31708]=37;
cos[31709]=37;
cos[31710]=37;
cos[31711]=37;
cos[31712]=37;
cos[31713]=37;
cos[31714]=37;
cos[31715]=37;
cos[31716]=37;
cos[31717]=37;
cos[31718]=37;
cos[31719]=37;
cos[31720]=37;
cos[31721]=37;
cos[31722]=37;
cos[31723]=37;
cos[31724]=37;
cos[31725]=37;
cos[31726]=37;
cos[31727]=36;
cos[31728]=36;
cos[31729]=36;
cos[31730]=36;
cos[31731]=36;
cos[31732]=36;
cos[31733]=36;
cos[31734]=36;
cos[31735]=36;
cos[31736]=36;
cos[31737]=36;
cos[31738]=36;
cos[31739]=36;
cos[31740]=36;
cos[31741]=36;
cos[31742]=36;
cos[31743]=36;
cos[31744]=36;
cos[31745]=36;
cos[31746]=36;
cos[31747]=36;
cos[31748]=36;
cos[31749]=36;
cos[31750]=35;
cos[31751]=35;
cos[31752]=35;
cos[31753]=35;
cos[31754]=35;
cos[31755]=35;
cos[31756]=35;
cos[31757]=35;
cos[31758]=35;
cos[31759]=35;
cos[31760]=35;
cos[31761]=35;
cos[31762]=35;
cos[31763]=35;
cos[31764]=35;
cos[31765]=35;
cos[31766]=35;
cos[31767]=35;
cos[31768]=35;
cos[31769]=35;
cos[31770]=35;
cos[31771]=35;
cos[31772]=35;
cos[31773]=34;
cos[31774]=34;
cos[31775]=34;
cos[31776]=34;
cos[31777]=34;
cos[31778]=34;
cos[31779]=34;
cos[31780]=34;
cos[31781]=34;
cos[31782]=34;
cos[31783]=34;
cos[31784]=34;
cos[31785]=34;
cos[31786]=34;
cos[31787]=34;
cos[31788]=34;
cos[31789]=34;
cos[31790]=34;
cos[31791]=34;
cos[31792]=34;
cos[31793]=34;
cos[31794]=34;
cos[31795]=33;
cos[31796]=33;
cos[31797]=33;
cos[31798]=33;
cos[31799]=33;
cos[31800]=33;
cos[31801]=33;
cos[31802]=33;
cos[31803]=33;
cos[31804]=33;
cos[31805]=33;
cos[31806]=33;
cos[31807]=33;
cos[31808]=33;
cos[31809]=33;
cos[31810]=33;
cos[31811]=33;
cos[31812]=33;
cos[31813]=33;
cos[31814]=33;
cos[31815]=33;
cos[31816]=33;
cos[31817]=33;
cos[31818]=32;
cos[31819]=32;
cos[31820]=32;
cos[31821]=32;
cos[31822]=32;
cos[31823]=32;
cos[31824]=32;
cos[31825]=32;
cos[31826]=32;
cos[31827]=32;
cos[31828]=32;
cos[31829]=32;
cos[31830]=32;
cos[31831]=32;
cos[31832]=32;
cos[31833]=32;
cos[31834]=32;
cos[31835]=32;
cos[31836]=32;
cos[31837]=32;
cos[31838]=32;
cos[31839]=32;
cos[31840]=31;
cos[31841]=31;
cos[31842]=31;
cos[31843]=31;
cos[31844]=31;
cos[31845]=31;
cos[31846]=31;
cos[31847]=31;
cos[31848]=31;
cos[31849]=31;
cos[31850]=31;
cos[31851]=31;
cos[31852]=31;
cos[31853]=31;
cos[31854]=31;
cos[31855]=31;
cos[31856]=31;
cos[31857]=31;
cos[31858]=31;
cos[31859]=31;
cos[31860]=31;
cos[31861]=31;
cos[31862]=30;
cos[31863]=30;
cos[31864]=30;
cos[31865]=30;
cos[31866]=30;
cos[31867]=30;
cos[31868]=30;
cos[31869]=30;
cos[31870]=30;
cos[31871]=30;
cos[31872]=30;
cos[31873]=30;
cos[31874]=30;
cos[31875]=30;
cos[31876]=30;
cos[31877]=30;
cos[31878]=30;
cos[31879]=30;
cos[31880]=30;
cos[31881]=30;
cos[31882]=30;
cos[31883]=30;
cos[31884]=29;
cos[31885]=29;
cos[31886]=29;
cos[31887]=29;
cos[31888]=29;
cos[31889]=29;
cos[31890]=29;
cos[31891]=29;
cos[31892]=29;
cos[31893]=29;
cos[31894]=29;
cos[31895]=29;
cos[31896]=29;
cos[31897]=29;
cos[31898]=29;
cos[31899]=29;
cos[31900]=29;
cos[31901]=29;
cos[31902]=29;
cos[31903]=29;
cos[31904]=29;
cos[31905]=29;
cos[31906]=28;
cos[31907]=28;
cos[31908]=28;
cos[31909]=28;
cos[31910]=28;
cos[31911]=28;
cos[31912]=28;
cos[31913]=28;
cos[31914]=28;
cos[31915]=28;
cos[31916]=28;
cos[31917]=28;
cos[31918]=28;
cos[31919]=28;
cos[31920]=28;
cos[31921]=28;
cos[31922]=28;
cos[31923]=28;
cos[31924]=28;
cos[31925]=28;
cos[31926]=28;
cos[31927]=28;
cos[31928]=27;
cos[31929]=27;
cos[31930]=27;
cos[31931]=27;
cos[31932]=27;
cos[31933]=27;
cos[31934]=27;
cos[31935]=27;
cos[31936]=27;
cos[31937]=27;
cos[31938]=27;
cos[31939]=27;
cos[31940]=27;
cos[31941]=27;
cos[31942]=27;
cos[31943]=27;
cos[31944]=27;
cos[31945]=27;
cos[31946]=27;
cos[31947]=27;
cos[31948]=27;
cos[31949]=27;
cos[31950]=26;
cos[31951]=26;
cos[31952]=26;
cos[31953]=26;
cos[31954]=26;
cos[31955]=26;
cos[31956]=26;
cos[31957]=26;
cos[31958]=26;
cos[31959]=26;
cos[31960]=26;
cos[31961]=26;
cos[31962]=26;
cos[31963]=26;
cos[31964]=26;
cos[31965]=26;
cos[31966]=26;
cos[31967]=26;
cos[31968]=26;
cos[31969]=26;
cos[31970]=26;
cos[31971]=25;
cos[31972]=25;
cos[31973]=25;
cos[31974]=25;
cos[31975]=25;
cos[31976]=25;
cos[31977]=25;
cos[31978]=25;
cos[31979]=25;
cos[31980]=25;
cos[31981]=25;
cos[31982]=25;
cos[31983]=25;
cos[31984]=25;
cos[31985]=25;
cos[31986]=25;
cos[31987]=25;
cos[31988]=25;
cos[31989]=25;
cos[31990]=25;
cos[31991]=25;
cos[31992]=25;
cos[31993]=24;
cos[31994]=24;
cos[31995]=24;
cos[31996]=24;
cos[31997]=24;
cos[31998]=24;
cos[31999]=24;
cos[32000]=24;
cos[32001]=24;
cos[32002]=24;
cos[32003]=24;
cos[32004]=24;
cos[32005]=24;
cos[32006]=24;
cos[32007]=24;
cos[32008]=24;
cos[32009]=24;
cos[32010]=24;
cos[32011]=24;
cos[32012]=24;
cos[32013]=24;
cos[32014]=23;
cos[32015]=23;
cos[32016]=23;
cos[32017]=23;
cos[32018]=23;
cos[32019]=23;
cos[32020]=23;
cos[32021]=23;
cos[32022]=23;
cos[32023]=23;
cos[32024]=23;
cos[32025]=23;
cos[32026]=23;
cos[32027]=23;
cos[32028]=23;
cos[32029]=23;
cos[32030]=23;
cos[32031]=23;
cos[32032]=23;
cos[32033]=23;
cos[32034]=23;
cos[32035]=23;
cos[32036]=22;
cos[32037]=22;
cos[32038]=22;
cos[32039]=22;
cos[32040]=22;
cos[32041]=22;
cos[32042]=22;
cos[32043]=22;
cos[32044]=22;
cos[32045]=22;
cos[32046]=22;
cos[32047]=22;
cos[32048]=22;
cos[32049]=22;
cos[32050]=22;
cos[32051]=22;
cos[32052]=22;
cos[32053]=22;
cos[32054]=22;
cos[32055]=22;
cos[32056]=22;
cos[32057]=21;
cos[32058]=21;
cos[32059]=21;
cos[32060]=21;
cos[32061]=21;
cos[32062]=21;
cos[32063]=21;
cos[32064]=21;
cos[32065]=21;
cos[32066]=21;
cos[32067]=21;
cos[32068]=21;
cos[32069]=21;
cos[32070]=21;
cos[32071]=21;
cos[32072]=21;
cos[32073]=21;
cos[32074]=21;
cos[32075]=21;
cos[32076]=21;
cos[32077]=21;
cos[32078]=20;
cos[32079]=20;
cos[32080]=20;
cos[32081]=20;
cos[32082]=20;
cos[32083]=20;
cos[32084]=20;
cos[32085]=20;
cos[32086]=20;
cos[32087]=20;
cos[32088]=20;
cos[32089]=20;
cos[32090]=20;
cos[32091]=20;
cos[32092]=20;
cos[32093]=20;
cos[32094]=20;
cos[32095]=20;
cos[32096]=20;
cos[32097]=20;
cos[32098]=20;
cos[32099]=19;
cos[32100]=19;
cos[32101]=19;
cos[32102]=19;
cos[32103]=19;
cos[32104]=19;
cos[32105]=19;
cos[32106]=19;
cos[32107]=19;
cos[32108]=19;
cos[32109]=19;
cos[32110]=19;
cos[32111]=19;
cos[32112]=19;
cos[32113]=19;
cos[32114]=19;
cos[32115]=19;
cos[32116]=19;
cos[32117]=19;
cos[32118]=19;
cos[32119]=19;
cos[32120]=18;
cos[32121]=18;
cos[32122]=18;
cos[32123]=18;
cos[32124]=18;
cos[32125]=18;
cos[32126]=18;
cos[32127]=18;
cos[32128]=18;
cos[32129]=18;
cos[32130]=18;
cos[32131]=18;
cos[32132]=18;
cos[32133]=18;
cos[32134]=18;
cos[32135]=18;
cos[32136]=18;
cos[32137]=18;
cos[32138]=18;
cos[32139]=18;
cos[32140]=18;
cos[32141]=17;
cos[32142]=17;
cos[32143]=17;
cos[32144]=17;
cos[32145]=17;
cos[32146]=17;
cos[32147]=17;
cos[32148]=17;
cos[32149]=17;
cos[32150]=17;
cos[32151]=17;
cos[32152]=17;
cos[32153]=17;
cos[32154]=17;
cos[32155]=17;
cos[32156]=17;
cos[32157]=17;
cos[32158]=17;
cos[32159]=17;
cos[32160]=17;
cos[32161]=17;
cos[32162]=16;
cos[32163]=16;
cos[32164]=16;
cos[32165]=16;
cos[32166]=16;
cos[32167]=16;
cos[32168]=16;
cos[32169]=16;
cos[32170]=16;
cos[32171]=16;
cos[32172]=16;
cos[32173]=16;
cos[32174]=16;
cos[32175]=16;
cos[32176]=16;
cos[32177]=16;
cos[32178]=16;
cos[32179]=16;
cos[32180]=16;
cos[32181]=16;
cos[32182]=16;
cos[32183]=15;
cos[32184]=15;
cos[32185]=15;
cos[32186]=15;
cos[32187]=15;
cos[32188]=15;
cos[32189]=15;
cos[32190]=15;
cos[32191]=15;
cos[32192]=15;
cos[32193]=15;
cos[32194]=15;
cos[32195]=15;
cos[32196]=15;
cos[32197]=15;
cos[32198]=15;
cos[32199]=15;
cos[32200]=15;
cos[32201]=15;
cos[32202]=15;
cos[32203]=14;
cos[32204]=14;
cos[32205]=14;
cos[32206]=14;
cos[32207]=14;
cos[32208]=14;
cos[32209]=14;
cos[32210]=14;
cos[32211]=14;
cos[32212]=14;
cos[32213]=14;
cos[32214]=14;
cos[32215]=14;
cos[32216]=14;
cos[32217]=14;
cos[32218]=14;
cos[32219]=14;
cos[32220]=14;
cos[32221]=14;
cos[32222]=14;
cos[32223]=14;
cos[32224]=13;
cos[32225]=13;
cos[32226]=13;
cos[32227]=13;
cos[32228]=13;
cos[32229]=13;
cos[32230]=13;
cos[32231]=13;
cos[32232]=13;
cos[32233]=13;
cos[32234]=13;
cos[32235]=13;
cos[32236]=13;
cos[32237]=13;
cos[32238]=13;
cos[32239]=13;
cos[32240]=13;
cos[32241]=13;
cos[32242]=13;
cos[32243]=13;
cos[32244]=13;
cos[32245]=12;
cos[32246]=12;
cos[32247]=12;
cos[32248]=12;
cos[32249]=12;
cos[32250]=12;
cos[32251]=12;
cos[32252]=12;
cos[32253]=12;
cos[32254]=12;
cos[32255]=12;
cos[32256]=12;
cos[32257]=12;
cos[32258]=12;
cos[32259]=12;
cos[32260]=12;
cos[32261]=12;
cos[32262]=12;
cos[32263]=12;
cos[32264]=12;
cos[32265]=11;
cos[32266]=11;
cos[32267]=11;
cos[32268]=11;
cos[32269]=11;
cos[32270]=11;
cos[32271]=11;
cos[32272]=11;
cos[32273]=11;
cos[32274]=11;
cos[32275]=11;
cos[32276]=11;
cos[32277]=11;
cos[32278]=11;
cos[32279]=11;
cos[32280]=11;
cos[32281]=11;
cos[32282]=11;
cos[32283]=11;
cos[32284]=11;
cos[32285]=11;
cos[32286]=10;
cos[32287]=10;
cos[32288]=10;
cos[32289]=10;
cos[32290]=10;
cos[32291]=10;
cos[32292]=10;
cos[32293]=10;
cos[32294]=10;
cos[32295]=10;
cos[32296]=10;
cos[32297]=10;
cos[32298]=10;
cos[32299]=10;
cos[32300]=10;
cos[32301]=10;
cos[32302]=10;
cos[32303]=10;
cos[32304]=10;
cos[32305]=10;
cos[32306]=9;
cos[32307]=9;
cos[32308]=9;
cos[32309]=9;
cos[32310]=9;
cos[32311]=9;
cos[32312]=9;
cos[32313]=9;
cos[32314]=9;
cos[32315]=9;
cos[32316]=9;
cos[32317]=9;
cos[32318]=9;
cos[32319]=9;
cos[32320]=9;
cos[32321]=9;
cos[32322]=9;
cos[32323]=9;
cos[32324]=9;
cos[32325]=9;
cos[32326]=9;
cos[32327]=8;
cos[32328]=8;
cos[32329]=8;
cos[32330]=8;
cos[32331]=8;
cos[32332]=8;
cos[32333]=8;
cos[32334]=8;
cos[32335]=8;
cos[32336]=8;
cos[32337]=8;
cos[32338]=8;
cos[32339]=8;
cos[32340]=8;
cos[32341]=8;
cos[32342]=8;
cos[32343]=8;
cos[32344]=8;
cos[32345]=8;
cos[32346]=8;
cos[32347]=7;
cos[32348]=7;
cos[32349]=7;
cos[32350]=7;
cos[32351]=7;
cos[32352]=7;
cos[32353]=7;
cos[32354]=7;
cos[32355]=7;
cos[32356]=7;
cos[32357]=7;
cos[32358]=7;
cos[32359]=7;
cos[32360]=7;
cos[32361]=7;
cos[32362]=7;
cos[32363]=7;
cos[32364]=7;
cos[32365]=7;
cos[32366]=7;
cos[32367]=7;
cos[32368]=6;
cos[32369]=6;
cos[32370]=6;
cos[32371]=6;
cos[32372]=6;
cos[32373]=6;
cos[32374]=6;
cos[32375]=6;
cos[32376]=6;
cos[32377]=6;
cos[32378]=6;
cos[32379]=6;
cos[32380]=6;
cos[32381]=6;
cos[32382]=6;
cos[32383]=6;
cos[32384]=6;
cos[32385]=6;
cos[32386]=6;
cos[32387]=6;
cos[32388]=5;
cos[32389]=5;
cos[32390]=5;
cos[32391]=5;
cos[32392]=5;
cos[32393]=5;
cos[32394]=5;
cos[32395]=5;
cos[32396]=5;
cos[32397]=5;
cos[32398]=5;
cos[32399]=5;
cos[32400]=5;
cos[32401]=5;
cos[32402]=5;
cos[32403]=5;
cos[32404]=5;
cos[32405]=5;
cos[32406]=5;
cos[32407]=5;
cos[32408]=5;
cos[32409]=4;
cos[32410]=4;
cos[32411]=4;
cos[32412]=4;
cos[32413]=4;
cos[32414]=4;
cos[32415]=4;
cos[32416]=4;
cos[32417]=4;
cos[32418]=4;
cos[32419]=4;
cos[32420]=4;
cos[32421]=4;
cos[32422]=4;
cos[32423]=4;
cos[32424]=4;
cos[32425]=4;
cos[32426]=4;
cos[32427]=4;
cos[32428]=4;
cos[32429]=3;
cos[32430]=3;
cos[32431]=3;
cos[32432]=3;
cos[32433]=3;
cos[32434]=3;
cos[32435]=3;
cos[32436]=3;
cos[32437]=3;
cos[32438]=3;
cos[32439]=3;
cos[32440]=3;
cos[32441]=3;
cos[32442]=3;
cos[32443]=3;
cos[32444]=3;
cos[32445]=3;
cos[32446]=3;
cos[32447]=3;
cos[32448]=3;
cos[32449]=3;
cos[32450]=2;
cos[32451]=2;
cos[32452]=2;
cos[32453]=2;
cos[32454]=2;
cos[32455]=2;
cos[32456]=2;
cos[32457]=2;
cos[32458]=2;
cos[32459]=2;
cos[32460]=2;
cos[32461]=2;
cos[32462]=2;
cos[32463]=2;
cos[32464]=2;
cos[32465]=2;
cos[32466]=2;
cos[32467]=2;
cos[32468]=2;
cos[32469]=2;
cos[32470]=1;
cos[32471]=1;
cos[32472]=1;
cos[32473]=1;
cos[32474]=1;
cos[32475]=1;
cos[32476]=1;
cos[32477]=1;
cos[32478]=1;
cos[32479]=1;
cos[32480]=1;
cos[32481]=1;
cos[32482]=1;
cos[32483]=1;
cos[32484]=1;
cos[32485]=1;
cos[32486]=1;
cos[32487]=1;
cos[32488]=1;
cos[32489]=1;
cos[32490]=0;
cos[32491]=0;
cos[32492]=0;
cos[32493]=0;
cos[32494]=0;
cos[32495]=0;
cos[32496]=0;
cos[32497]=0;
cos[32498]=0;
cos[32499]=0;
cos[32500]=0;
cos[32501]=0;
cos[32502]=0;
cos[32503]=0;
cos[32504]=0;
cos[32505]=0;
cos[32506]=0;
cos[32507]=0;
cos[32508]=0;
cos[32509]=0;
cos[32510]=0;
cos[32511]=-1;
cos[32512]=-1;
cos[32513]=-1;
cos[32514]=-1;
cos[32515]=-1;
cos[32516]=-1;
cos[32517]=-1;
cos[32518]=-1;
cos[32519]=-1;
cos[32520]=-1;
cos[32521]=-1;
cos[32522]=-1;
cos[32523]=-1;
cos[32524]=-1;
cos[32525]=-1;
cos[32526]=-1;
cos[32527]=-1;
cos[32528]=-1;
cos[32529]=-1;
cos[32530]=-1;
cos[32531]=-2;
cos[32532]=-2;
cos[32533]=-2;
cos[32534]=-2;
cos[32535]=-2;
cos[32536]=-2;
cos[32537]=-2;
cos[32538]=-2;
cos[32539]=-2;
cos[32540]=-2;
cos[32541]=-2;
cos[32542]=-2;
cos[32543]=-2;
cos[32544]=-2;
cos[32545]=-2;
cos[32546]=-2;
cos[32547]=-2;
cos[32548]=-2;
cos[32549]=-2;
cos[32550]=-2;
cos[32551]=-3;
cos[32552]=-3;
cos[32553]=-3;
cos[32554]=-3;
cos[32555]=-3;
cos[32556]=-3;
cos[32557]=-3;
cos[32558]=-3;
cos[32559]=-3;
cos[32560]=-3;
cos[32561]=-3;
cos[32562]=-3;
cos[32563]=-3;
cos[32564]=-3;
cos[32565]=-3;
cos[32566]=-3;
cos[32567]=-3;
cos[32568]=-3;
cos[32569]=-3;
cos[32570]=-3;
cos[32571]=-3;
cos[32572]=-4;
cos[32573]=-4;
cos[32574]=-4;
cos[32575]=-4;
cos[32576]=-4;
cos[32577]=-4;
cos[32578]=-4;
cos[32579]=-4;
cos[32580]=-4;
cos[32581]=-4;
cos[32582]=-4;
cos[32583]=-4;
cos[32584]=-4;
cos[32585]=-4;
cos[32586]=-4;
cos[32587]=-4;
cos[32588]=-4;
cos[32589]=-4;
cos[32590]=-4;
cos[32591]=-4;
cos[32592]=-5;
cos[32593]=-5;
cos[32594]=-5;
cos[32595]=-5;
cos[32596]=-5;
cos[32597]=-5;
cos[32598]=-5;
cos[32599]=-5;
cos[32600]=-5;
cos[32601]=-5;
cos[32602]=-5;
cos[32603]=-5;
cos[32604]=-5;
cos[32605]=-5;
cos[32606]=-5;
cos[32607]=-5;
cos[32608]=-5;
cos[32609]=-5;
cos[32610]=-5;
cos[32611]=-5;
cos[32612]=-5;
cos[32613]=-6;
cos[32614]=-6;
cos[32615]=-6;
cos[32616]=-6;
cos[32617]=-6;
cos[32618]=-6;
cos[32619]=-6;
cos[32620]=-6;
cos[32621]=-6;
cos[32622]=-6;
cos[32623]=-6;
cos[32624]=-6;
cos[32625]=-6;
cos[32626]=-6;
cos[32627]=-6;
cos[32628]=-6;
cos[32629]=-6;
cos[32630]=-6;
cos[32631]=-6;
cos[32632]=-6;
cos[32633]=-7;
cos[32634]=-7;
cos[32635]=-7;
cos[32636]=-7;
cos[32637]=-7;
cos[32638]=-7;
cos[32639]=-7;
cos[32640]=-7;
cos[32641]=-7;
cos[32642]=-7;
cos[32643]=-7;
cos[32644]=-7;
cos[32645]=-7;
cos[32646]=-7;
cos[32647]=-7;
cos[32648]=-7;
cos[32649]=-7;
cos[32650]=-7;
cos[32651]=-7;
cos[32652]=-7;
cos[32653]=-7;
cos[32654]=-8;
cos[32655]=-8;
cos[32656]=-8;
cos[32657]=-8;
cos[32658]=-8;
cos[32659]=-8;
cos[32660]=-8;
cos[32661]=-8;
cos[32662]=-8;
cos[32663]=-8;
cos[32664]=-8;
cos[32665]=-8;
cos[32666]=-8;
cos[32667]=-8;
cos[32668]=-8;
cos[32669]=-8;
cos[32670]=-8;
cos[32671]=-8;
cos[32672]=-8;
cos[32673]=-8;
cos[32674]=-9;
cos[32675]=-9;
cos[32676]=-9;
cos[32677]=-9;
cos[32678]=-9;
cos[32679]=-9;
cos[32680]=-9;
cos[32681]=-9;
cos[32682]=-9;
cos[32683]=-9;
cos[32684]=-9;
cos[32685]=-9;
cos[32686]=-9;
cos[32687]=-9;
cos[32688]=-9;
cos[32689]=-9;
cos[32690]=-9;
cos[32691]=-9;
cos[32692]=-9;
cos[32693]=-9;
cos[32694]=-9;
cos[32695]=-10;
cos[32696]=-10;
cos[32697]=-10;
cos[32698]=-10;
cos[32699]=-10;
cos[32700]=-10;
cos[32701]=-10;
cos[32702]=-10;
cos[32703]=-10;
cos[32704]=-10;
cos[32705]=-10;
cos[32706]=-10;
cos[32707]=-10;
cos[32708]=-10;
cos[32709]=-10;
cos[32710]=-10;
cos[32711]=-10;
cos[32712]=-10;
cos[32713]=-10;
cos[32714]=-10;
cos[32715]=-11;
cos[32716]=-11;
cos[32717]=-11;
cos[32718]=-11;
cos[32719]=-11;
cos[32720]=-11;
cos[32721]=-11;
cos[32722]=-11;
cos[32723]=-11;
cos[32724]=-11;
cos[32725]=-11;
cos[32726]=-11;
cos[32727]=-11;
cos[32728]=-11;
cos[32729]=-11;
cos[32730]=-11;
cos[32731]=-11;
cos[32732]=-11;
cos[32733]=-11;
cos[32734]=-11;
cos[32735]=-11;
cos[32736]=-12;
cos[32737]=-12;
cos[32738]=-12;
cos[32739]=-12;
cos[32740]=-12;
cos[32741]=-12;
cos[32742]=-12;
cos[32743]=-12;
cos[32744]=-12;
cos[32745]=-12;
cos[32746]=-12;
cos[32747]=-12;
cos[32748]=-12;
cos[32749]=-12;
cos[32750]=-12;
cos[32751]=-12;
cos[32752]=-12;
cos[32753]=-12;
cos[32754]=-12;
cos[32755]=-12;
cos[32756]=-13;
cos[32757]=-13;
cos[32758]=-13;
cos[32759]=-13;
cos[32760]=-13;
cos[32761]=-13;
cos[32762]=-13;
cos[32763]=-13;
cos[32764]=-13;
cos[32765]=-13;
cos[32766]=-13;
cos[32767]=-13;
cos[32768]=-13;
cos[32769]=-13;
cos[32770]=-13;
cos[32771]=-13;
cos[32772]=-13;
cos[32773]=-13;
cos[32774]=-13;
cos[32775]=-13;
cos[32776]=-13;
cos[32777]=-14;
cos[32778]=-14;
cos[32779]=-14;
cos[32780]=-14;
cos[32781]=-14;
cos[32782]=-14;
cos[32783]=-14;
cos[32784]=-14;
cos[32785]=-14;
cos[32786]=-14;
cos[32787]=-14;
cos[32788]=-14;
cos[32789]=-14;
cos[32790]=-14;
cos[32791]=-14;
cos[32792]=-14;
cos[32793]=-14;
cos[32794]=-14;
cos[32795]=-14;
cos[32796]=-14;
cos[32797]=-14;
cos[32798]=-15;
cos[32799]=-15;
cos[32800]=-15;
cos[32801]=-15;
cos[32802]=-15;
cos[32803]=-15;
cos[32804]=-15;
cos[32805]=-15;
cos[32806]=-15;
cos[32807]=-15;
cos[32808]=-15;
cos[32809]=-15;
cos[32810]=-15;
cos[32811]=-15;
cos[32812]=-15;
cos[32813]=-15;
cos[32814]=-15;
cos[32815]=-15;
cos[32816]=-15;
cos[32817]=-15;
cos[32818]=-16;
cos[32819]=-16;
cos[32820]=-16;
cos[32821]=-16;
cos[32822]=-16;
cos[32823]=-16;
cos[32824]=-16;
cos[32825]=-16;
cos[32826]=-16;
cos[32827]=-16;
cos[32828]=-16;
cos[32829]=-16;
cos[32830]=-16;
cos[32831]=-16;
cos[32832]=-16;
cos[32833]=-16;
cos[32834]=-16;
cos[32835]=-16;
cos[32836]=-16;
cos[32837]=-16;
cos[32838]=-16;
cos[32839]=-17;
cos[32840]=-17;
cos[32841]=-17;
cos[32842]=-17;
cos[32843]=-17;
cos[32844]=-17;
cos[32845]=-17;
cos[32846]=-17;
cos[32847]=-17;
cos[32848]=-17;
cos[32849]=-17;
cos[32850]=-17;
cos[32851]=-17;
cos[32852]=-17;
cos[32853]=-17;
cos[32854]=-17;
cos[32855]=-17;
cos[32856]=-17;
cos[32857]=-17;
cos[32858]=-17;
cos[32859]=-17;
cos[32860]=-18;
cos[32861]=-18;
cos[32862]=-18;
cos[32863]=-18;
cos[32864]=-18;
cos[32865]=-18;
cos[32866]=-18;
cos[32867]=-18;
cos[32868]=-18;
cos[32869]=-18;
cos[32870]=-18;
cos[32871]=-18;
cos[32872]=-18;
cos[32873]=-18;
cos[32874]=-18;
cos[32875]=-18;
cos[32876]=-18;
cos[32877]=-18;
cos[32878]=-18;
cos[32879]=-18;
cos[32880]=-18;
cos[32881]=-19;
cos[32882]=-19;
cos[32883]=-19;
cos[32884]=-19;
cos[32885]=-19;
cos[32886]=-19;
cos[32887]=-19;
cos[32888]=-19;
cos[32889]=-19;
cos[32890]=-19;
cos[32891]=-19;
cos[32892]=-19;
cos[32893]=-19;
cos[32894]=-19;
cos[32895]=-19;
cos[32896]=-19;
cos[32897]=-19;
cos[32898]=-19;
cos[32899]=-19;
cos[32900]=-19;
cos[32901]=-19;
cos[32902]=-20;
cos[32903]=-20;
cos[32904]=-20;
cos[32905]=-20;
cos[32906]=-20;
cos[32907]=-20;
cos[32908]=-20;
cos[32909]=-20;
cos[32910]=-20;
cos[32911]=-20;
cos[32912]=-20;
cos[32913]=-20;
cos[32914]=-20;
cos[32915]=-20;
cos[32916]=-20;
cos[32917]=-20;
cos[32918]=-20;
cos[32919]=-20;
cos[32920]=-20;
cos[32921]=-20;
cos[32922]=-20;
cos[32923]=-21;
cos[32924]=-21;
cos[32925]=-21;
cos[32926]=-21;
cos[32927]=-21;
cos[32928]=-21;
cos[32929]=-21;
cos[32930]=-21;
cos[32931]=-21;
cos[32932]=-21;
cos[32933]=-21;
cos[32934]=-21;
cos[32935]=-21;
cos[32936]=-21;
cos[32937]=-21;
cos[32938]=-21;
cos[32939]=-21;
cos[32940]=-21;
cos[32941]=-21;
cos[32942]=-21;
cos[32943]=-21;
cos[32944]=-22;
cos[32945]=-22;
cos[32946]=-22;
cos[32947]=-22;
cos[32948]=-22;
cos[32949]=-22;
cos[32950]=-22;
cos[32951]=-22;
cos[32952]=-22;
cos[32953]=-22;
cos[32954]=-22;
cos[32955]=-22;
cos[32956]=-22;
cos[32957]=-22;
cos[32958]=-22;
cos[32959]=-22;
cos[32960]=-22;
cos[32961]=-22;
cos[32962]=-22;
cos[32963]=-22;
cos[32964]=-22;
cos[32965]=-23;
cos[32966]=-23;
cos[32967]=-23;
cos[32968]=-23;
cos[32969]=-23;
cos[32970]=-23;
cos[32971]=-23;
cos[32972]=-23;
cos[32973]=-23;
cos[32974]=-23;
cos[32975]=-23;
cos[32976]=-23;
cos[32977]=-23;
cos[32978]=-23;
cos[32979]=-23;
cos[32980]=-23;
cos[32981]=-23;
cos[32982]=-23;
cos[32983]=-23;
cos[32984]=-23;
cos[32985]=-23;
cos[32986]=-23;
cos[32987]=-24;
cos[32988]=-24;
cos[32989]=-24;
cos[32990]=-24;
cos[32991]=-24;
cos[32992]=-24;
cos[32993]=-24;
cos[32994]=-24;
cos[32995]=-24;
cos[32996]=-24;
cos[32997]=-24;
cos[32998]=-24;
cos[32999]=-24;
cos[33000]=-24;
cos[33001]=-24;
cos[33002]=-24;
cos[33003]=-24;
cos[33004]=-24;
cos[33005]=-24;
cos[33006]=-24;
cos[33007]=-24;
cos[33008]=-25;
cos[33009]=-25;
cos[33010]=-25;
cos[33011]=-25;
cos[33012]=-25;
cos[33013]=-25;
cos[33014]=-25;
cos[33015]=-25;
cos[33016]=-25;
cos[33017]=-25;
cos[33018]=-25;
cos[33019]=-25;
cos[33020]=-25;
cos[33021]=-25;
cos[33022]=-25;
cos[33023]=-25;
cos[33024]=-25;
cos[33025]=-25;
cos[33026]=-25;
cos[33027]=-25;
cos[33028]=-25;
cos[33029]=-25;
cos[33030]=-26;
cos[33031]=-26;
cos[33032]=-26;
cos[33033]=-26;
cos[33034]=-26;
cos[33035]=-26;
cos[33036]=-26;
cos[33037]=-26;
cos[33038]=-26;
cos[33039]=-26;
cos[33040]=-26;
cos[33041]=-26;
cos[33042]=-26;
cos[33043]=-26;
cos[33044]=-26;
cos[33045]=-26;
cos[33046]=-26;
cos[33047]=-26;
cos[33048]=-26;
cos[33049]=-26;
cos[33050]=-26;
cos[33051]=-27;
cos[33052]=-27;
cos[33053]=-27;
cos[33054]=-27;
cos[33055]=-27;
cos[33056]=-27;
cos[33057]=-27;
cos[33058]=-27;
cos[33059]=-27;
cos[33060]=-27;
cos[33061]=-27;
cos[33062]=-27;
cos[33063]=-27;
cos[33064]=-27;
cos[33065]=-27;
cos[33066]=-27;
cos[33067]=-27;
cos[33068]=-27;
cos[33069]=-27;
cos[33070]=-27;
cos[33071]=-27;
cos[33072]=-27;
cos[33073]=-28;
cos[33074]=-28;
cos[33075]=-28;
cos[33076]=-28;
cos[33077]=-28;
cos[33078]=-28;
cos[33079]=-28;
cos[33080]=-28;
cos[33081]=-28;
cos[33082]=-28;
cos[33083]=-28;
cos[33084]=-28;
cos[33085]=-28;
cos[33086]=-28;
cos[33087]=-28;
cos[33088]=-28;
cos[33089]=-28;
cos[33090]=-28;
cos[33091]=-28;
cos[33092]=-28;
cos[33093]=-28;
cos[33094]=-28;
cos[33095]=-29;
cos[33096]=-29;
cos[33097]=-29;
cos[33098]=-29;
cos[33099]=-29;
cos[33100]=-29;
cos[33101]=-29;
cos[33102]=-29;
cos[33103]=-29;
cos[33104]=-29;
cos[33105]=-29;
cos[33106]=-29;
cos[33107]=-29;
cos[33108]=-29;
cos[33109]=-29;
cos[33110]=-29;
cos[33111]=-29;
cos[33112]=-29;
cos[33113]=-29;
cos[33114]=-29;
cos[33115]=-29;
cos[33116]=-29;
cos[33117]=-30;
cos[33118]=-30;
cos[33119]=-30;
cos[33120]=-30;
cos[33121]=-30;
cos[33122]=-30;
cos[33123]=-30;
cos[33124]=-30;
cos[33125]=-30;
cos[33126]=-30;
cos[33127]=-30;
cos[33128]=-30;
cos[33129]=-30;
cos[33130]=-30;
cos[33131]=-30;
cos[33132]=-30;
cos[33133]=-30;
cos[33134]=-30;
cos[33135]=-30;
cos[33136]=-30;
cos[33137]=-30;
cos[33138]=-30;
cos[33139]=-31;
cos[33140]=-31;
cos[33141]=-31;
cos[33142]=-31;
cos[33143]=-31;
cos[33144]=-31;
cos[33145]=-31;
cos[33146]=-31;
cos[33147]=-31;
cos[33148]=-31;
cos[33149]=-31;
cos[33150]=-31;
cos[33151]=-31;
cos[33152]=-31;
cos[33153]=-31;
cos[33154]=-31;
cos[33155]=-31;
cos[33156]=-31;
cos[33157]=-31;
cos[33158]=-31;
cos[33159]=-31;
cos[33160]=-31;
cos[33161]=-32;
cos[33162]=-32;
cos[33163]=-32;
cos[33164]=-32;
cos[33165]=-32;
cos[33166]=-32;
cos[33167]=-32;
cos[33168]=-32;
cos[33169]=-32;
cos[33170]=-32;
cos[33171]=-32;
cos[33172]=-32;
cos[33173]=-32;
cos[33174]=-32;
cos[33175]=-32;
cos[33176]=-32;
cos[33177]=-32;
cos[33178]=-32;
cos[33179]=-32;
cos[33180]=-32;
cos[33181]=-32;
cos[33182]=-32;
cos[33183]=-33;
cos[33184]=-33;
cos[33185]=-33;
cos[33186]=-33;
cos[33187]=-33;
cos[33188]=-33;
cos[33189]=-33;
cos[33190]=-33;
cos[33191]=-33;
cos[33192]=-33;
cos[33193]=-33;
cos[33194]=-33;
cos[33195]=-33;
cos[33196]=-33;
cos[33197]=-33;
cos[33198]=-33;
cos[33199]=-33;
cos[33200]=-33;
cos[33201]=-33;
cos[33202]=-33;
cos[33203]=-33;
cos[33204]=-33;
cos[33205]=-33;
cos[33206]=-34;
cos[33207]=-34;
cos[33208]=-34;
cos[33209]=-34;
cos[33210]=-34;
cos[33211]=-34;
cos[33212]=-34;
cos[33213]=-34;
cos[33214]=-34;
cos[33215]=-34;
cos[33216]=-34;
cos[33217]=-34;
cos[33218]=-34;
cos[33219]=-34;
cos[33220]=-34;
cos[33221]=-34;
cos[33222]=-34;
cos[33223]=-34;
cos[33224]=-34;
cos[33225]=-34;
cos[33226]=-34;
cos[33227]=-34;
cos[33228]=-35;
cos[33229]=-35;
cos[33230]=-35;
cos[33231]=-35;
cos[33232]=-35;
cos[33233]=-35;
cos[33234]=-35;
cos[33235]=-35;
cos[33236]=-35;
cos[33237]=-35;
cos[33238]=-35;
cos[33239]=-35;
cos[33240]=-35;
cos[33241]=-35;
cos[33242]=-35;
cos[33243]=-35;
cos[33244]=-35;
cos[33245]=-35;
cos[33246]=-35;
cos[33247]=-35;
cos[33248]=-35;
cos[33249]=-35;
cos[33250]=-35;
cos[33251]=-36;
cos[33252]=-36;
cos[33253]=-36;
cos[33254]=-36;
cos[33255]=-36;
cos[33256]=-36;
cos[33257]=-36;
cos[33258]=-36;
cos[33259]=-36;
cos[33260]=-36;
cos[33261]=-36;
cos[33262]=-36;
cos[33263]=-36;
cos[33264]=-36;
cos[33265]=-36;
cos[33266]=-36;
cos[33267]=-36;
cos[33268]=-36;
cos[33269]=-36;
cos[33270]=-36;
cos[33271]=-36;
cos[33272]=-36;
cos[33273]=-36;
cos[33274]=-37;
cos[33275]=-37;
cos[33276]=-37;
cos[33277]=-37;
cos[33278]=-37;
cos[33279]=-37;
cos[33280]=-37;
cos[33281]=-37;
cos[33282]=-37;
cos[33283]=-37;
cos[33284]=-37;
cos[33285]=-37;
cos[33286]=-37;
cos[33287]=-37;
cos[33288]=-37;
cos[33289]=-37;
cos[33290]=-37;
cos[33291]=-37;
cos[33292]=-37;
cos[33293]=-37;
cos[33294]=-37;
cos[33295]=-37;
cos[33296]=-37;
cos[33297]=-38;
cos[33298]=-38;
cos[33299]=-38;
cos[33300]=-38;
cos[33301]=-38;
cos[33302]=-38;
cos[33303]=-38;
cos[33304]=-38;
cos[33305]=-38;
cos[33306]=-38;
cos[33307]=-38;
cos[33308]=-38;
cos[33309]=-38;
cos[33310]=-38;
cos[33311]=-38;
cos[33312]=-38;
cos[33313]=-38;
cos[33314]=-38;
cos[33315]=-38;
cos[33316]=-38;
cos[33317]=-38;
cos[33318]=-38;
cos[33319]=-38;
cos[33320]=-38;
cos[33321]=-39;
cos[33322]=-39;
cos[33323]=-39;
cos[33324]=-39;
cos[33325]=-39;
cos[33326]=-39;
cos[33327]=-39;
cos[33328]=-39;
cos[33329]=-39;
cos[33330]=-39;
cos[33331]=-39;
cos[33332]=-39;
cos[33333]=-39;
cos[33334]=-39;
cos[33335]=-39;
cos[33336]=-39;
cos[33337]=-39;
cos[33338]=-39;
cos[33339]=-39;
cos[33340]=-39;
cos[33341]=-39;
cos[33342]=-39;
cos[33343]=-39;
cos[33344]=-40;
cos[33345]=-40;
cos[33346]=-40;
cos[33347]=-40;
cos[33348]=-40;
cos[33349]=-40;
cos[33350]=-40;
cos[33351]=-40;
cos[33352]=-40;
cos[33353]=-40;
cos[33354]=-40;
cos[33355]=-40;
cos[33356]=-40;
cos[33357]=-40;
cos[33358]=-40;
cos[33359]=-40;
cos[33360]=-40;
cos[33361]=-40;
cos[33362]=-40;
cos[33363]=-40;
cos[33364]=-40;
cos[33365]=-40;
cos[33366]=-40;
cos[33367]=-40;
cos[33368]=-41;
cos[33369]=-41;
cos[33370]=-41;
cos[33371]=-41;
cos[33372]=-41;
cos[33373]=-41;
cos[33374]=-41;
cos[33375]=-41;
cos[33376]=-41;
cos[33377]=-41;
cos[33378]=-41;
cos[33379]=-41;
cos[33380]=-41;
cos[33381]=-41;
cos[33382]=-41;
cos[33383]=-41;
cos[33384]=-41;
cos[33385]=-41;
cos[33386]=-41;
cos[33387]=-41;
cos[33388]=-41;
cos[33389]=-41;
cos[33390]=-41;
cos[33391]=-41;
cos[33392]=-42;
cos[33393]=-42;
cos[33394]=-42;
cos[33395]=-42;
cos[33396]=-42;
cos[33397]=-42;
cos[33398]=-42;
cos[33399]=-42;
cos[33400]=-42;
cos[33401]=-42;
cos[33402]=-42;
cos[33403]=-42;
cos[33404]=-42;
cos[33405]=-42;
cos[33406]=-42;
cos[33407]=-42;
cos[33408]=-42;
cos[33409]=-42;
cos[33410]=-42;
cos[33411]=-42;
cos[33412]=-42;
cos[33413]=-42;
cos[33414]=-42;
cos[33415]=-42;
cos[33416]=-43;
cos[33417]=-43;
cos[33418]=-43;
cos[33419]=-43;
cos[33420]=-43;
cos[33421]=-43;
cos[33422]=-43;
cos[33423]=-43;
cos[33424]=-43;
cos[33425]=-43;
cos[33426]=-43;
cos[33427]=-43;
cos[33428]=-43;
cos[33429]=-43;
cos[33430]=-43;
cos[33431]=-43;
cos[33432]=-43;
cos[33433]=-43;
cos[33434]=-43;
cos[33435]=-43;
cos[33436]=-43;
cos[33437]=-43;
cos[33438]=-43;
cos[33439]=-43;
cos[33440]=-44;
cos[33441]=-44;
cos[33442]=-44;
cos[33443]=-44;
cos[33444]=-44;
cos[33445]=-44;
cos[33446]=-44;
cos[33447]=-44;
cos[33448]=-44;
cos[33449]=-44;
cos[33450]=-44;
cos[33451]=-44;
cos[33452]=-44;
cos[33453]=-44;
cos[33454]=-44;
cos[33455]=-44;
cos[33456]=-44;
cos[33457]=-44;
cos[33458]=-44;
cos[33459]=-44;
cos[33460]=-44;
cos[33461]=-44;
cos[33462]=-44;
cos[33463]=-44;
cos[33464]=-44;
cos[33465]=-45;
cos[33466]=-45;
cos[33467]=-45;
cos[33468]=-45;
cos[33469]=-45;
cos[33470]=-45;
cos[33471]=-45;
cos[33472]=-45;
cos[33473]=-45;
cos[33474]=-45;
cos[33475]=-45;
cos[33476]=-45;
cos[33477]=-45;
cos[33478]=-45;
cos[33479]=-45;
cos[33480]=-45;
cos[33481]=-45;
cos[33482]=-45;
cos[33483]=-45;
cos[33484]=-45;
cos[33485]=-45;
cos[33486]=-45;
cos[33487]=-45;
cos[33488]=-45;
cos[33489]=-45;
cos[33490]=-46;
cos[33491]=-46;
cos[33492]=-46;
cos[33493]=-46;
cos[33494]=-46;
cos[33495]=-46;
cos[33496]=-46;
cos[33497]=-46;
cos[33498]=-46;
cos[33499]=-46;
cos[33500]=-46;
cos[33501]=-46;
cos[33502]=-46;
cos[33503]=-46;
cos[33504]=-46;
cos[33505]=-46;
cos[33506]=-46;
cos[33507]=-46;
cos[33508]=-46;
cos[33509]=-46;
cos[33510]=-46;
cos[33511]=-46;
cos[33512]=-46;
cos[33513]=-46;
cos[33514]=-46;
cos[33515]=-47;
cos[33516]=-47;
cos[33517]=-47;
cos[33518]=-47;
cos[33519]=-47;
cos[33520]=-47;
cos[33521]=-47;
cos[33522]=-47;
cos[33523]=-47;
cos[33524]=-47;
cos[33525]=-47;
cos[33526]=-47;
cos[33527]=-47;
cos[33528]=-47;
cos[33529]=-47;
cos[33530]=-47;
cos[33531]=-47;
cos[33532]=-47;
cos[33533]=-47;
cos[33534]=-47;
cos[33535]=-47;
cos[33536]=-47;
cos[33537]=-47;
cos[33538]=-47;
cos[33539]=-47;
cos[33540]=-47;
cos[33541]=-48;
cos[33542]=-48;
cos[33543]=-48;
cos[33544]=-48;
cos[33545]=-48;
cos[33546]=-48;
cos[33547]=-48;
cos[33548]=-48;
cos[33549]=-48;
cos[33550]=-48;
cos[33551]=-48;
cos[33552]=-48;
cos[33553]=-48;
cos[33554]=-48;
cos[33555]=-48;
cos[33556]=-48;
cos[33557]=-48;
cos[33558]=-48;
cos[33559]=-48;
cos[33560]=-48;
cos[33561]=-48;
cos[33562]=-48;
cos[33563]=-48;
cos[33564]=-48;
cos[33565]=-48;
cos[33566]=-49;
cos[33567]=-49;
cos[33568]=-49;
cos[33569]=-49;
cos[33570]=-49;
cos[33571]=-49;
cos[33572]=-49;
cos[33573]=-49;
cos[33574]=-49;
cos[33575]=-49;
cos[33576]=-49;
cos[33577]=-49;
cos[33578]=-49;
cos[33579]=-49;
cos[33580]=-49;
cos[33581]=-49;
cos[33582]=-49;
cos[33583]=-49;
cos[33584]=-49;
cos[33585]=-49;
cos[33586]=-49;
cos[33587]=-49;
cos[33588]=-49;
cos[33589]=-49;
cos[33590]=-49;
cos[33591]=-49;
cos[33592]=-49;
cos[33593]=-50;
cos[33594]=-50;
cos[33595]=-50;
cos[33596]=-50;
cos[33597]=-50;
cos[33598]=-50;
cos[33599]=-50;
cos[33600]=-50;
cos[33601]=-50;
cos[33602]=-50;
cos[33603]=-50;
cos[33604]=-50;
cos[33605]=-50;
cos[33606]=-50;
cos[33607]=-50;
cos[33608]=-50;
cos[33609]=-50;
cos[33610]=-50;
cos[33611]=-50;
cos[33612]=-50;
cos[33613]=-50;
cos[33614]=-50;
cos[33615]=-50;
cos[33616]=-50;
cos[33617]=-50;
cos[33618]=-50;
cos[33619]=-51;
cos[33620]=-51;
cos[33621]=-51;
cos[33622]=-51;
cos[33623]=-51;
cos[33624]=-51;
cos[33625]=-51;
cos[33626]=-51;
cos[33627]=-51;
cos[33628]=-51;
cos[33629]=-51;
cos[33630]=-51;
cos[33631]=-51;
cos[33632]=-51;
cos[33633]=-51;
cos[33634]=-51;
cos[33635]=-51;
cos[33636]=-51;
cos[33637]=-51;
cos[33638]=-51;
cos[33639]=-51;
cos[33640]=-51;
cos[33641]=-51;
cos[33642]=-51;
cos[33643]=-51;
cos[33644]=-51;
cos[33645]=-51;
cos[33646]=-52;
cos[33647]=-52;
cos[33648]=-52;
cos[33649]=-52;
cos[33650]=-52;
cos[33651]=-52;
cos[33652]=-52;
cos[33653]=-52;
cos[33654]=-52;
cos[33655]=-52;
cos[33656]=-52;
cos[33657]=-52;
cos[33658]=-52;
cos[33659]=-52;
cos[33660]=-52;
cos[33661]=-52;
cos[33662]=-52;
cos[33663]=-52;
cos[33664]=-52;
cos[33665]=-52;
cos[33666]=-52;
cos[33667]=-52;
cos[33668]=-52;
cos[33669]=-52;
cos[33670]=-52;
cos[33671]=-52;
cos[33672]=-52;
cos[33673]=-53;
cos[33674]=-53;
cos[33675]=-53;
cos[33676]=-53;
cos[33677]=-53;
cos[33678]=-53;
cos[33679]=-53;
cos[33680]=-53;
cos[33681]=-53;
cos[33682]=-53;
cos[33683]=-53;
cos[33684]=-53;
cos[33685]=-53;
cos[33686]=-53;
cos[33687]=-53;
cos[33688]=-53;
cos[33689]=-53;
cos[33690]=-53;
cos[33691]=-53;
cos[33692]=-53;
cos[33693]=-53;
cos[33694]=-53;
cos[33695]=-53;
cos[33696]=-53;
cos[33697]=-53;
cos[33698]=-53;
cos[33699]=-53;
cos[33700]=-53;
cos[33701]=-54;
cos[33702]=-54;
cos[33703]=-54;
cos[33704]=-54;
cos[33705]=-54;
cos[33706]=-54;
cos[33707]=-54;
cos[33708]=-54;
cos[33709]=-54;
cos[33710]=-54;
cos[33711]=-54;
cos[33712]=-54;
cos[33713]=-54;
cos[33714]=-54;
cos[33715]=-54;
cos[33716]=-54;
cos[33717]=-54;
cos[33718]=-54;
cos[33719]=-54;
cos[33720]=-54;
cos[33721]=-54;
cos[33722]=-54;
cos[33723]=-54;
cos[33724]=-54;
cos[33725]=-54;
cos[33726]=-54;
cos[33727]=-54;
cos[33728]=-54;
cos[33729]=-55;
cos[33730]=-55;
cos[33731]=-55;
cos[33732]=-55;
cos[33733]=-55;
cos[33734]=-55;
cos[33735]=-55;
cos[33736]=-55;
cos[33737]=-55;
cos[33738]=-55;
cos[33739]=-55;
cos[33740]=-55;
cos[33741]=-55;
cos[33742]=-55;
cos[33743]=-55;
cos[33744]=-55;
cos[33745]=-55;
cos[33746]=-55;
cos[33747]=-55;
cos[33748]=-55;
cos[33749]=-55;
cos[33750]=-55;
cos[33751]=-55;
cos[33752]=-55;
cos[33753]=-55;
cos[33754]=-55;
cos[33755]=-55;
cos[33756]=-55;
cos[33757]=-55;
cos[33758]=-56;
cos[33759]=-56;
cos[33760]=-56;
cos[33761]=-56;
cos[33762]=-56;
cos[33763]=-56;
cos[33764]=-56;
cos[33765]=-56;
cos[33766]=-56;
cos[33767]=-56;
cos[33768]=-56;
cos[33769]=-56;
cos[33770]=-56;
cos[33771]=-56;
cos[33772]=-56;
cos[33773]=-56;
cos[33774]=-56;
cos[33775]=-56;
cos[33776]=-56;
cos[33777]=-56;
cos[33778]=-56;
cos[33779]=-56;
cos[33780]=-56;
cos[33781]=-56;
cos[33782]=-56;
cos[33783]=-56;
cos[33784]=-56;
cos[33785]=-56;
cos[33786]=-56;
cos[33787]=-57;
cos[33788]=-57;
cos[33789]=-57;
cos[33790]=-57;
cos[33791]=-57;
cos[33792]=-57;
cos[33793]=-57;
cos[33794]=-57;
cos[33795]=-57;
cos[33796]=-57;
cos[33797]=-57;
cos[33798]=-57;
cos[33799]=-57;
cos[33800]=-57;
cos[33801]=-57;
cos[33802]=-57;
cos[33803]=-57;
cos[33804]=-57;
cos[33805]=-57;
cos[33806]=-57;
cos[33807]=-57;
cos[33808]=-57;
cos[33809]=-57;
cos[33810]=-57;
cos[33811]=-57;
cos[33812]=-57;
cos[33813]=-57;
cos[33814]=-57;
cos[33815]=-57;
cos[33816]=-57;
cos[33817]=-58;
cos[33818]=-58;
cos[33819]=-58;
cos[33820]=-58;
cos[33821]=-58;
cos[33822]=-58;
cos[33823]=-58;
cos[33824]=-58;
cos[33825]=-58;
cos[33826]=-58;
cos[33827]=-58;
cos[33828]=-58;
cos[33829]=-58;
cos[33830]=-58;
cos[33831]=-58;
cos[33832]=-58;
cos[33833]=-58;
cos[33834]=-58;
cos[33835]=-58;
cos[33836]=-58;
cos[33837]=-58;
cos[33838]=-58;
cos[33839]=-58;
cos[33840]=-58;
cos[33841]=-58;
cos[33842]=-58;
cos[33843]=-58;
cos[33844]=-58;
cos[33845]=-58;
cos[33846]=-58;
cos[33847]=-59;
cos[33848]=-59;
cos[33849]=-59;
cos[33850]=-59;
cos[33851]=-59;
cos[33852]=-59;
cos[33853]=-59;
cos[33854]=-59;
cos[33855]=-59;
cos[33856]=-59;
cos[33857]=-59;
cos[33858]=-59;
cos[33859]=-59;
cos[33860]=-59;
cos[33861]=-59;
cos[33862]=-59;
cos[33863]=-59;
cos[33864]=-59;
cos[33865]=-59;
cos[33866]=-59;
cos[33867]=-59;
cos[33868]=-59;
cos[33869]=-59;
cos[33870]=-59;
cos[33871]=-59;
cos[33872]=-59;
cos[33873]=-59;
cos[33874]=-59;
cos[33875]=-59;
cos[33876]=-59;
cos[33877]=-59;
cos[33878]=-60;
cos[33879]=-60;
cos[33880]=-60;
cos[33881]=-60;
cos[33882]=-60;
cos[33883]=-60;
cos[33884]=-60;
cos[33885]=-60;
cos[33886]=-60;
cos[33887]=-60;
cos[33888]=-60;
cos[33889]=-60;
cos[33890]=-60;
cos[33891]=-60;
cos[33892]=-60;
cos[33893]=-60;
cos[33894]=-60;
cos[33895]=-60;
cos[33896]=-60;
cos[33897]=-60;
cos[33898]=-60;
cos[33899]=-60;
cos[33900]=-60;
cos[33901]=-60;
cos[33902]=-60;
cos[33903]=-60;
cos[33904]=-60;
cos[33905]=-60;
cos[33906]=-60;
cos[33907]=-60;
cos[33908]=-60;
cos[33909]=-60;
cos[33910]=-61;
cos[33911]=-61;
cos[33912]=-61;
cos[33913]=-61;
cos[33914]=-61;
cos[33915]=-61;
cos[33916]=-61;
cos[33917]=-61;
cos[33918]=-61;
cos[33919]=-61;
cos[33920]=-61;
cos[33921]=-61;
cos[33922]=-61;
cos[33923]=-61;
cos[33924]=-61;
cos[33925]=-61;
cos[33926]=-61;
cos[33927]=-61;
cos[33928]=-61;
cos[33929]=-61;
cos[33930]=-61;
cos[33931]=-61;
cos[33932]=-61;
cos[33933]=-61;
cos[33934]=-61;
cos[33935]=-61;
cos[33936]=-61;
cos[33937]=-61;
cos[33938]=-61;
cos[33939]=-61;
cos[33940]=-61;
cos[33941]=-61;
cos[33942]=-61;
cos[33943]=-62;
cos[33944]=-62;
cos[33945]=-62;
cos[33946]=-62;
cos[33947]=-62;
cos[33948]=-62;
cos[33949]=-62;
cos[33950]=-62;
cos[33951]=-62;
cos[33952]=-62;
cos[33953]=-62;
cos[33954]=-62;
cos[33955]=-62;
cos[33956]=-62;
cos[33957]=-62;
cos[33958]=-62;
cos[33959]=-62;
cos[33960]=-62;
cos[33961]=-62;
cos[33962]=-62;
cos[33963]=-62;
cos[33964]=-62;
cos[33965]=-62;
cos[33966]=-62;
cos[33967]=-62;
cos[33968]=-62;
cos[33969]=-62;
cos[33970]=-62;
cos[33971]=-62;
cos[33972]=-62;
cos[33973]=-62;
cos[33974]=-62;
cos[33975]=-62;
cos[33976]=-63;
cos[33977]=-63;
cos[33978]=-63;
cos[33979]=-63;
cos[33980]=-63;
cos[33981]=-63;
cos[33982]=-63;
cos[33983]=-63;
cos[33984]=-63;
cos[33985]=-63;
cos[33986]=-63;
cos[33987]=-63;
cos[33988]=-63;
cos[33989]=-63;
cos[33990]=-63;
cos[33991]=-63;
cos[33992]=-63;
cos[33993]=-63;
cos[33994]=-63;
cos[33995]=-63;
cos[33996]=-63;
cos[33997]=-63;
cos[33998]=-63;
cos[33999]=-63;
cos[34000]=-63;
cos[34001]=-63;
cos[34002]=-63;
cos[34003]=-63;
cos[34004]=-63;
cos[34005]=-63;
cos[34006]=-63;
cos[34007]=-63;
cos[34008]=-63;
cos[34009]=-63;
cos[34010]=-63;
cos[34011]=-64;
cos[34012]=-64;
cos[34013]=-64;
cos[34014]=-64;
cos[34015]=-64;
cos[34016]=-64;
cos[34017]=-64;
cos[34018]=-64;
cos[34019]=-64;
cos[34020]=-64;
cos[34021]=-64;
cos[34022]=-64;
cos[34023]=-64;
cos[34024]=-64;
cos[34025]=-64;
cos[34026]=-64;
cos[34027]=-64;
cos[34028]=-64;
cos[34029]=-64;
cos[34030]=-64;
cos[34031]=-64;
cos[34032]=-64;
cos[34033]=-64;
cos[34034]=-64;
cos[34035]=-64;
cos[34036]=-64;
cos[34037]=-64;
cos[34038]=-64;
cos[34039]=-64;
cos[34040]=-64;
cos[34041]=-64;
cos[34042]=-64;
cos[34043]=-64;
cos[34044]=-64;
cos[34045]=-64;
cos[34046]=-65;
cos[34047]=-65;
cos[34048]=-65;
cos[34049]=-65;
cos[34050]=-65;
cos[34051]=-65;
cos[34052]=-65;
cos[34053]=-65;
cos[34054]=-65;
cos[34055]=-65;
cos[34056]=-65;
cos[34057]=-65;
cos[34058]=-65;
cos[34059]=-65;
cos[34060]=-65;
cos[34061]=-65;
cos[34062]=-65;
cos[34063]=-65;
cos[34064]=-65;
cos[34065]=-65;
cos[34066]=-65;
cos[34067]=-65;
cos[34068]=-65;
cos[34069]=-65;
cos[34070]=-65;
cos[34071]=-65;
cos[34072]=-65;
cos[34073]=-65;
cos[34074]=-65;
cos[34075]=-65;
cos[34076]=-65;
cos[34077]=-65;
cos[34078]=-65;
cos[34079]=-65;
cos[34080]=-65;
cos[34081]=-65;
cos[34082]=-65;
cos[34083]=-66;
cos[34084]=-66;
cos[34085]=-66;
cos[34086]=-66;
cos[34087]=-66;
cos[34088]=-66;
cos[34089]=-66;
cos[34090]=-66;
cos[34091]=-66;
cos[34092]=-66;
cos[34093]=-66;
cos[34094]=-66;
cos[34095]=-66;
cos[34096]=-66;
cos[34097]=-66;
cos[34098]=-66;
cos[34099]=-66;
cos[34100]=-66;
cos[34101]=-66;
cos[34102]=-66;
cos[34103]=-66;
cos[34104]=-66;
cos[34105]=-66;
cos[34106]=-66;
cos[34107]=-66;
cos[34108]=-66;
cos[34109]=-66;
cos[34110]=-66;
cos[34111]=-66;
cos[34112]=-66;
cos[34113]=-66;
cos[34114]=-66;
cos[34115]=-66;
cos[34116]=-66;
cos[34117]=-66;
cos[34118]=-66;
cos[34119]=-66;
cos[34120]=-66;
cos[34121]=-67;
cos[34122]=-67;
cos[34123]=-67;
cos[34124]=-67;
cos[34125]=-67;
cos[34126]=-67;
cos[34127]=-67;
cos[34128]=-67;
cos[34129]=-67;
cos[34130]=-67;
cos[34131]=-67;
cos[34132]=-67;
cos[34133]=-67;
cos[34134]=-67;
cos[34135]=-67;
cos[34136]=-67;
cos[34137]=-67;
cos[34138]=-67;
cos[34139]=-67;
cos[34140]=-67;
cos[34141]=-67;
cos[34142]=-67;
cos[34143]=-67;
cos[34144]=-67;
cos[34145]=-67;
cos[34146]=-67;
cos[34147]=-67;
cos[34148]=-67;
cos[34149]=-67;
cos[34150]=-67;
cos[34151]=-67;
cos[34152]=-67;
cos[34153]=-67;
cos[34154]=-67;
cos[34155]=-67;
cos[34156]=-67;
cos[34157]=-67;
cos[34158]=-67;
cos[34159]=-67;
cos[34160]=-67;
cos[34161]=-68;
cos[34162]=-68;
cos[34163]=-68;
cos[34164]=-68;
cos[34165]=-68;
cos[34166]=-68;
cos[34167]=-68;
cos[34168]=-68;
cos[34169]=-68;
cos[34170]=-68;
cos[34171]=-68;
cos[34172]=-68;
cos[34173]=-68;
cos[34174]=-68;
cos[34175]=-68;
cos[34176]=-68;
cos[34177]=-68;
cos[34178]=-68;
cos[34179]=-68;
cos[34180]=-68;
cos[34181]=-68;
cos[34182]=-68;
cos[34183]=-68;
cos[34184]=-68;
cos[34185]=-68;
cos[34186]=-68;
cos[34187]=-68;
cos[34188]=-68;
cos[34189]=-68;
cos[34190]=-68;
cos[34191]=-68;
cos[34192]=-68;
cos[34193]=-68;
cos[34194]=-68;
cos[34195]=-68;
cos[34196]=-68;
cos[34197]=-68;
cos[34198]=-68;
cos[34199]=-68;
cos[34200]=-68;
cos[34201]=-68;
cos[34202]=-69;
cos[34203]=-69;
cos[34204]=-69;
cos[34205]=-69;
cos[34206]=-69;
cos[34207]=-69;
cos[34208]=-69;
cos[34209]=-69;
cos[34210]=-69;
cos[34211]=-69;
cos[34212]=-69;
cos[34213]=-69;
cos[34214]=-69;
cos[34215]=-69;
cos[34216]=-69;
cos[34217]=-69;
cos[34218]=-69;
cos[34219]=-69;
cos[34220]=-69;
cos[34221]=-69;
cos[34222]=-69;
cos[34223]=-69;
cos[34224]=-69;
cos[34225]=-69;
cos[34226]=-69;
cos[34227]=-69;
cos[34228]=-69;
cos[34229]=-69;
cos[34230]=-69;
cos[34231]=-69;
cos[34232]=-69;
cos[34233]=-69;
cos[34234]=-69;
cos[34235]=-69;
cos[34236]=-69;
cos[34237]=-69;
cos[34238]=-69;
cos[34239]=-69;
cos[34240]=-69;
cos[34241]=-69;
cos[34242]=-69;
cos[34243]=-69;
cos[34244]=-69;
cos[34245]=-69;
cos[34246]=-70;
cos[34247]=-70;
cos[34248]=-70;
cos[34249]=-70;
cos[34250]=-70;
cos[34251]=-70;
cos[34252]=-70;
cos[34253]=-70;
cos[34254]=-70;
cos[34255]=-70;
cos[34256]=-70;
cos[34257]=-70;
cos[34258]=-70;
cos[34259]=-70;
cos[34260]=-70;
cos[34261]=-70;
cos[34262]=-70;
cos[34263]=-70;
cos[34264]=-70;
cos[34265]=-70;
cos[34266]=-70;
cos[34267]=-70;
cos[34268]=-70;
cos[34269]=-70;
cos[34270]=-70;
cos[34271]=-70;
cos[34272]=-70;
cos[34273]=-70;
cos[34274]=-70;
cos[34275]=-70;
cos[34276]=-70;
cos[34277]=-70;
cos[34278]=-70;
cos[34279]=-70;
cos[34280]=-70;
cos[34281]=-70;
cos[34282]=-70;
cos[34283]=-70;
cos[34284]=-70;
cos[34285]=-70;
cos[34286]=-70;
cos[34287]=-70;
cos[34288]=-70;
cos[34289]=-70;
cos[34290]=-70;
cos[34291]=-71;
cos[34292]=-71;
cos[34293]=-71;
cos[34294]=-71;
cos[34295]=-71;
cos[34296]=-71;
cos[34297]=-71;
cos[34298]=-71;
cos[34299]=-71;
cos[34300]=-71;
cos[34301]=-71;
cos[34302]=-71;
cos[34303]=-71;
cos[34304]=-71;
cos[34305]=-71;
cos[34306]=-71;
cos[34307]=-71;
cos[34308]=-71;
cos[34309]=-71;
cos[34310]=-71;
cos[34311]=-71;
cos[34312]=-71;
cos[34313]=-71;
cos[34314]=-71;
cos[34315]=-71;
cos[34316]=-71;
cos[34317]=-71;
cos[34318]=-71;
cos[34319]=-71;
cos[34320]=-71;
cos[34321]=-71;
cos[34322]=-71;
cos[34323]=-71;
cos[34324]=-71;
cos[34325]=-71;
cos[34326]=-71;
cos[34327]=-71;
cos[34328]=-71;
cos[34329]=-71;
cos[34330]=-71;
cos[34331]=-71;
cos[34332]=-71;
cos[34333]=-71;
cos[34334]=-71;
cos[34335]=-71;
cos[34336]=-71;
cos[34337]=-71;
cos[34338]=-71;
cos[34339]=-71;
cos[34340]=-72;
cos[34341]=-72;
cos[34342]=-72;
cos[34343]=-72;
cos[34344]=-72;
cos[34345]=-72;
cos[34346]=-72;
cos[34347]=-72;
cos[34348]=-72;
cos[34349]=-72;
cos[34350]=-72;
cos[34351]=-72;
cos[34352]=-72;
cos[34353]=-72;
cos[34354]=-72;
cos[34355]=-72;
cos[34356]=-72;
cos[34357]=-72;
cos[34358]=-72;
cos[34359]=-72;
cos[34360]=-72;
cos[34361]=-72;
cos[34362]=-72;
cos[34363]=-72;
cos[34364]=-72;
cos[34365]=-72;
cos[34366]=-72;
cos[34367]=-72;
cos[34368]=-72;
cos[34369]=-72;
cos[34370]=-72;
cos[34371]=-72;
cos[34372]=-72;
cos[34373]=-72;
cos[34374]=-72;
cos[34375]=-72;
cos[34376]=-72;
cos[34377]=-72;
cos[34378]=-72;
cos[34379]=-72;
cos[34380]=-72;
cos[34381]=-72;
cos[34382]=-72;
cos[34383]=-72;
cos[34384]=-72;
cos[34385]=-72;
cos[34386]=-72;
cos[34387]=-72;
cos[34388]=-72;
cos[34389]=-72;
cos[34390]=-72;
cos[34391]=-72;
cos[34392]=-72;
cos[34393]=-73;
cos[34394]=-73;
cos[34395]=-73;
cos[34396]=-73;
cos[34397]=-73;
cos[34398]=-73;
cos[34399]=-73;
cos[34400]=-73;
cos[34401]=-73;
cos[34402]=-73;
cos[34403]=-73;
cos[34404]=-73;
cos[34405]=-73;
cos[34406]=-73;
cos[34407]=-73;
cos[34408]=-73;
cos[34409]=-73;
cos[34410]=-73;
cos[34411]=-73;
cos[34412]=-73;
cos[34413]=-73;
cos[34414]=-73;
cos[34415]=-73;
cos[34416]=-73;
cos[34417]=-73;
cos[34418]=-73;
cos[34419]=-73;
cos[34420]=-73;
cos[34421]=-73;
cos[34422]=-73;
cos[34423]=-73;
cos[34424]=-73;
cos[34425]=-73;
cos[34426]=-73;
cos[34427]=-73;
cos[34428]=-73;
cos[34429]=-73;
cos[34430]=-73;
cos[34431]=-73;
cos[34432]=-73;
cos[34433]=-73;
cos[34434]=-73;
cos[34435]=-73;
cos[34436]=-73;
cos[34437]=-73;
cos[34438]=-73;
cos[34439]=-73;
cos[34440]=-73;
cos[34441]=-73;
cos[34442]=-73;
cos[34443]=-73;
cos[34444]=-73;
cos[34445]=-73;
cos[34446]=-73;
cos[34447]=-73;
cos[34448]=-73;
cos[34449]=-73;
cos[34450]=-74;
cos[34451]=-74;
cos[34452]=-74;
cos[34453]=-74;
cos[34454]=-74;
cos[34455]=-74;
cos[34456]=-74;
cos[34457]=-74;
cos[34458]=-74;
cos[34459]=-74;
cos[34460]=-74;
cos[34461]=-74;
cos[34462]=-74;
cos[34463]=-74;
cos[34464]=-74;
cos[34465]=-74;
cos[34466]=-74;
cos[34467]=-74;
cos[34468]=-74;
cos[34469]=-74;
cos[34470]=-74;
cos[34471]=-74;
cos[34472]=-74;
cos[34473]=-74;
cos[34474]=-74;
cos[34475]=-74;
cos[34476]=-74;
cos[34477]=-74;
cos[34478]=-74;
cos[34479]=-74;
cos[34480]=-74;
cos[34481]=-74;
cos[34482]=-74;
cos[34483]=-74;
cos[34484]=-74;
cos[34485]=-74;
cos[34486]=-74;
cos[34487]=-74;
cos[34488]=-74;
cos[34489]=-74;
cos[34490]=-74;
cos[34491]=-74;
cos[34492]=-74;
cos[34493]=-74;
cos[34494]=-74;
cos[34495]=-74;
cos[34496]=-74;
cos[34497]=-74;
cos[34498]=-74;
cos[34499]=-74;
cos[34500]=-74;
cos[34501]=-74;
cos[34502]=-74;
cos[34503]=-74;
cos[34504]=-74;
cos[34505]=-74;
cos[34506]=-74;
cos[34507]=-74;
cos[34508]=-74;
cos[34509]=-74;
cos[34510]=-74;
cos[34511]=-74;
cos[34512]=-74;
cos[34513]=-74;
cos[34514]=-75;
cos[34515]=-75;
cos[34516]=-75;
cos[34517]=-75;
cos[34518]=-75;
cos[34519]=-75;
cos[34520]=-75;
cos[34521]=-75;
cos[34522]=-75;
cos[34523]=-75;
cos[34524]=-75;
cos[34525]=-75;
cos[34526]=-75;
cos[34527]=-75;
cos[34528]=-75;
cos[34529]=-75;
cos[34530]=-75;
cos[34531]=-75;
cos[34532]=-75;
cos[34533]=-75;
cos[34534]=-75;
cos[34535]=-75;
cos[34536]=-75;
cos[34537]=-75;
cos[34538]=-75;
cos[34539]=-75;
cos[34540]=-75;
cos[34541]=-75;
cos[34542]=-75;
cos[34543]=-75;
cos[34544]=-75;
cos[34545]=-75;
cos[34546]=-75;
cos[34547]=-75;
cos[34548]=-75;
cos[34549]=-75;
cos[34550]=-75;
cos[34551]=-75;
cos[34552]=-75;
cos[34553]=-75;
cos[34554]=-75;
cos[34555]=-75;
cos[34556]=-75;
cos[34557]=-75;
cos[34558]=-75;
cos[34559]=-75;
cos[34560]=-75;
cos[34561]=-75;
cos[34562]=-75;
cos[34563]=-75;
cos[34564]=-75;
cos[34565]=-75;
cos[34566]=-75;
cos[34567]=-75;
cos[34568]=-75;
cos[34569]=-75;
cos[34570]=-75;
cos[34571]=-75;
cos[34572]=-75;
cos[34573]=-75;
cos[34574]=-75;
cos[34575]=-75;
cos[34576]=-75;
cos[34577]=-75;
cos[34578]=-75;
cos[34579]=-75;
cos[34580]=-75;
cos[34581]=-75;
cos[34582]=-75;
cos[34583]=-75;
cos[34584]=-75;
cos[34585]=-75;
cos[34586]=-75;
cos[34587]=-76;
cos[34588]=-76;
cos[34589]=-76;
cos[34590]=-76;
cos[34591]=-76;
cos[34592]=-76;
cos[34593]=-76;
cos[34594]=-76;
cos[34595]=-76;
cos[34596]=-76;
cos[34597]=-76;
cos[34598]=-76;
cos[34599]=-76;
cos[34600]=-76;
cos[34601]=-76;
cos[34602]=-76;
cos[34603]=-76;
cos[34604]=-76;
cos[34605]=-76;
cos[34606]=-76;
cos[34607]=-76;
cos[34608]=-76;
cos[34609]=-76;
cos[34610]=-76;
cos[34611]=-76;
cos[34612]=-76;
cos[34613]=-76;
cos[34614]=-76;
cos[34615]=-76;
cos[34616]=-76;
cos[34617]=-76;
cos[34618]=-76;
cos[34619]=-76;
cos[34620]=-76;
cos[34621]=-76;
cos[34622]=-76;
cos[34623]=-76;
cos[34624]=-76;
cos[34625]=-76;
cos[34626]=-76;
cos[34627]=-76;
cos[34628]=-76;
cos[34629]=-76;
cos[34630]=-76;
cos[34631]=-76;
cos[34632]=-76;
cos[34633]=-76;
cos[34634]=-76;
cos[34635]=-76;
cos[34636]=-76;
cos[34637]=-76;
cos[34638]=-76;
cos[34639]=-76;
cos[34640]=-76;
cos[34641]=-76;
cos[34642]=-76;
cos[34643]=-76;
cos[34644]=-76;
cos[34645]=-76;
cos[34646]=-76;
cos[34647]=-76;
cos[34648]=-76;
cos[34649]=-76;
cos[34650]=-76;
cos[34651]=-76;
cos[34652]=-76;
cos[34653]=-76;
cos[34654]=-76;
cos[34655]=-76;
cos[34656]=-76;
cos[34657]=-76;
cos[34658]=-76;
cos[34659]=-76;
cos[34660]=-76;
cos[34661]=-76;
cos[34662]=-76;
cos[34663]=-76;
cos[34664]=-76;
cos[34665]=-76;
cos[34666]=-76;
cos[34667]=-76;
cos[34668]=-76;
cos[34669]=-76;
cos[34670]=-76;
cos[34671]=-76;
cos[34672]=-76;
cos[34673]=-76;
cos[34674]=-76;
cos[34675]=-77;
cos[34676]=-77;
cos[34677]=-77;
cos[34678]=-77;
cos[34679]=-77;
cos[34680]=-77;
cos[34681]=-77;
cos[34682]=-77;
cos[34683]=-77;
cos[34684]=-77;
cos[34685]=-77;
cos[34686]=-77;
cos[34687]=-77;
cos[34688]=-77;
cos[34689]=-77;
cos[34690]=-77;
cos[34691]=-77;
cos[34692]=-77;
cos[34693]=-77;
cos[34694]=-77;
cos[34695]=-77;
cos[34696]=-77;
cos[34697]=-77;
cos[34698]=-77;
cos[34699]=-77;
cos[34700]=-77;
cos[34701]=-77;
cos[34702]=-77;
cos[34703]=-77;
cos[34704]=-77;
cos[34705]=-77;
cos[34706]=-77;
cos[34707]=-77;
cos[34708]=-77;
cos[34709]=-77;
cos[34710]=-77;
cos[34711]=-77;
cos[34712]=-77;
cos[34713]=-77;
cos[34714]=-77;
cos[34715]=-77;
cos[34716]=-77;
cos[34717]=-77;
cos[34718]=-77;
cos[34719]=-77;
cos[34720]=-77;
cos[34721]=-77;
cos[34722]=-77;
cos[34723]=-77;
cos[34724]=-77;
cos[34725]=-77;
cos[34726]=-77;
cos[34727]=-77;
cos[34728]=-77;
cos[34729]=-77;
cos[34730]=-77;
cos[34731]=-77;
cos[34732]=-77;
cos[34733]=-77;
cos[34734]=-77;
cos[34735]=-77;
cos[34736]=-77;
cos[34737]=-77;
cos[34738]=-77;
cos[34739]=-77;
cos[34740]=-77;
cos[34741]=-77;
cos[34742]=-77;
cos[34743]=-77;
cos[34744]=-77;
cos[34745]=-77;
cos[34746]=-77;
cos[34747]=-77;
cos[34748]=-77;
cos[34749]=-77;
cos[34750]=-77;
cos[34751]=-77;
cos[34752]=-77;
cos[34753]=-77;
cos[34754]=-77;
cos[34755]=-77;
cos[34756]=-77;
cos[34757]=-77;
cos[34758]=-77;
cos[34759]=-77;
cos[34760]=-77;
cos[34761]=-77;
cos[34762]=-77;
cos[34763]=-77;
cos[34764]=-77;
cos[34765]=-77;
cos[34766]=-77;
cos[34767]=-77;
cos[34768]=-77;
cos[34769]=-77;
cos[34770]=-77;
cos[34771]=-77;
cos[34772]=-77;
cos[34773]=-77;
cos[34774]=-77;
cos[34775]=-77;
cos[34776]=-77;
cos[34777]=-77;
cos[34778]=-77;
cos[34779]=-77;
cos[34780]=-77;
cos[34781]=-77;
cos[34782]=-77;
cos[34783]=-77;
cos[34784]=-77;
cos[34785]=-77;
cos[34786]=-77;
cos[34787]=-77;
cos[34788]=-77;
cos[34789]=-77;
cos[34790]=-77;
cos[34791]=-77;
cos[34792]=-77;
cos[34793]=-77;
cos[34794]=-77;
cos[34795]=-77;
cos[34796]=-77;
cos[34797]=-77;
cos[34798]=-77;
cos[34799]=-78;
cos[34800]=-78;
cos[34801]=-78;
cos[34802]=-78;
cos[34803]=-78;
cos[34804]=-78;
cos[34805]=-78;
cos[34806]=-78;
cos[34807]=-78;
cos[34808]=-78;
cos[34809]=-78;
cos[34810]=-78;
cos[34811]=-78;
cos[34812]=-78;
cos[34813]=-78;
cos[34814]=-78;
cos[34815]=-78;
cos[34816]=-78;
cos[34817]=-78;
cos[34818]=-78;
cos[34819]=-78;
cos[34820]=-78;
cos[34821]=-78;
cos[34822]=-78;
cos[34823]=-78;
cos[34824]=-78;
cos[34825]=-78;
cos[34826]=-78;
cos[34827]=-78;
cos[34828]=-78;
cos[34829]=-78;
cos[34830]=-78;
cos[34831]=-78;
cos[34832]=-78;
cos[34833]=-78;
cos[34834]=-78;
cos[34835]=-78;
cos[34836]=-78;
cos[34837]=-78;
cos[34838]=-78;
cos[34839]=-78;
cos[34840]=-78;
cos[34841]=-78;
cos[34842]=-78;
cos[34843]=-78;
cos[34844]=-78;
cos[34845]=-78;
cos[34846]=-78;
cos[34847]=-78;
cos[34848]=-78;
cos[34849]=-78;
cos[34850]=-78;
cos[34851]=-78;
cos[34852]=-78;
cos[34853]=-78;
cos[34854]=-78;
cos[34855]=-78;
cos[34856]=-78;
cos[34857]=-78;
cos[34858]=-78;
cos[34859]=-78;
cos[34860]=-78;
cos[34861]=-78;
cos[34862]=-78;
cos[34863]=-78;
cos[34864]=-78;
cos[34865]=-78;
cos[34866]=-78;
cos[34867]=-78;
cos[34868]=-78;
cos[34869]=-78;
cos[34870]=-78;
cos[34871]=-78;
cos[34872]=-78;
cos[34873]=-78;
cos[34874]=-78;
cos[34875]=-78;
cos[34876]=-78;
cos[34877]=-78;
cos[34878]=-78;
cos[34879]=-78;
cos[34880]=-78;
cos[34881]=-78;
cos[34882]=-78;
cos[34883]=-78;
cos[34884]=-78;
cos[34885]=-78;
cos[34886]=-78;
cos[34887]=-78;
cos[34888]=-78;
cos[34889]=-78;
cos[34890]=-78;
cos[34891]=-78;
cos[34892]=-78;
cos[34893]=-78;
cos[34894]=-78;
cos[34895]=-78;
cos[34896]=-78;
cos[34897]=-78;
cos[34898]=-78;
cos[34899]=-78;
cos[34900]=-78;
cos[34901]=-78;
cos[34902]=-78;
cos[34903]=-78;
cos[34904]=-78;
cos[34905]=-78;
cos[34906]=-78;
cos[34907]=-78;
cos[34908]=-78;
cos[34909]=-78;
cos[34910]=-78;
cos[34911]=-78;
cos[34912]=-78;
cos[34913]=-78;
cos[34914]=-78;
cos[34915]=-78;
cos[34916]=-78;
cos[34917]=-78;
cos[34918]=-78;
cos[34919]=-78;
cos[34920]=-78;
cos[34921]=-78;
cos[34922]=-78;
cos[34923]=-78;
cos[34924]=-78;
cos[34925]=-78;
cos[34926]=-78;
cos[34927]=-78;
cos[34928]=-78;
cos[34929]=-78;
cos[34930]=-78;
cos[34931]=-78;
cos[34932]=-78;
cos[34933]=-78;
cos[34934]=-78;
cos[34935]=-78;
cos[34936]=-78;
cos[34937]=-78;
cos[34938]=-78;
cos[34939]=-78;
cos[34940]=-78;
cos[34941]=-78;
cos[34942]=-78;
cos[34943]=-78;
cos[34944]=-78;
cos[34945]=-78;
cos[34946]=-78;
cos[34947]=-78;
cos[34948]=-78;
cos[34949]=-78;
cos[34950]=-78;
cos[34951]=-78;
cos[34952]=-78;
cos[34953]=-78;
cos[34954]=-78;
cos[34955]=-78;
cos[34956]=-78;
cos[34957]=-78;
cos[34958]=-78;
cos[34959]=-78;
cos[34960]=-78;
cos[34961]=-78;
cos[34962]=-78;
cos[34963]=-78;
cos[34964]=-78;
cos[34965]=-78;
cos[34966]=-78;
cos[34967]=-78;
cos[34968]=-78;
cos[34969]=-78;
cos[34970]=-78;
cos[34971]=-78;
cos[34972]=-78;
cos[34973]=-78;
cos[34974]=-78;
cos[34975]=-78;
cos[34976]=-78;
cos[34977]=-78;
cos[34978]=-78;
cos[34979]=-78;
cos[34980]=-78;
cos[34981]=-78;
cos[34982]=-78;
cos[34983]=-78;
cos[34984]=-78;
cos[34985]=-78;
cos[34986]=-78;
cos[34987]=-78;
cos[34988]=-78;
cos[34989]=-78;
cos[34990]=-78;
cos[34991]=-78;
cos[34992]=-78;
cos[34993]=-78;
cos[34994]=-78;
cos[34995]=-78;
cos[34996]=-78;
cos[34997]=-78;
cos[34998]=-78;
cos[34999]=-78;
cos[35000]=-78;
cos[35001]=-78;
cos[35002]=-78;
cos[35003]=-78;
cos[35004]=-78;
cos[35005]=-78;
cos[35006]=-78;
cos[35007]=-78;
cos[35008]=-78;
cos[35009]=-78;
cos[35010]=-78;
cos[35011]=-78;
cos[35012]=-78;
cos[35013]=-78;
cos[35014]=-78;
cos[35015]=-78;
cos[35016]=-78;
cos[35017]=-78;
cos[35018]=-78;
cos[35019]=-78;
cos[35020]=-78;
cos[35021]=-78;
cos[35022]=-78;
cos[35023]=-78;
cos[35024]=-78;
cos[35025]=-78;
cos[35026]=-78;
cos[35027]=-78;
cos[35028]=-78;
cos[35029]=-78;
cos[35030]=-78;
cos[35031]=-78;
cos[35032]=-78;
cos[35033]=-78;
cos[35034]=-78;
cos[35035]=-78;
cos[35036]=-78;
cos[35037]=-78;
cos[35038]=-78;
cos[35039]=-78;
cos[35040]=-78;
cos[35041]=-78;
cos[35042]=-78;
cos[35043]=-78;
cos[35044]=-78;
cos[35045]=-78;
cos[35046]=-78;
cos[35047]=-78;
cos[35048]=-78;
cos[35049]=-78;
cos[35050]=-78;
cos[35051]=-78;
cos[35052]=-78;
cos[35053]=-78;
cos[35054]=-78;
cos[35055]=-78;
cos[35056]=-78;
cos[35057]=-78;
cos[35058]=-78;
cos[35059]=-78;
cos[35060]=-78;
cos[35061]=-78;
cos[35062]=-78;
cos[35063]=-78;
cos[35064]=-78;
cos[35065]=-78;
cos[35066]=-78;
cos[35067]=-78;
cos[35068]=-78;
cos[35069]=-78;
cos[35070]=-78;
cos[35071]=-78;
cos[35072]=-78;
cos[35073]=-78;
cos[35074]=-78;
cos[35075]=-78;
cos[35076]=-78;
cos[35077]=-78;
cos[35078]=-78;
cos[35079]=-78;
cos[35080]=-78;
cos[35081]=-78;
cos[35082]=-78;
cos[35083]=-78;
cos[35084]=-78;
cos[35085]=-78;
cos[35086]=-78;
cos[35087]=-78;
cos[35088]=-78;
cos[35089]=-78;
cos[35090]=-78;
cos[35091]=-78;
cos[35092]=-78;
cos[35093]=-78;
cos[35094]=-78;
cos[35095]=-78;
cos[35096]=-78;
cos[35097]=-78;
cos[35098]=-78;
cos[35099]=-78;
cos[35100]=-78;
cos[35101]=-78;
cos[35102]=-78;
cos[35103]=-78;
cos[35104]=-78;
cos[35105]=-78;
cos[35106]=-78;
cos[35107]=-78;
cos[35108]=-78;
cos[35109]=-78;
cos[35110]=-78;
cos[35111]=-78;
cos[35112]=-78;
cos[35113]=-78;
cos[35114]=-78;
cos[35115]=-78;
cos[35116]=-78;
cos[35117]=-78;
cos[35118]=-78;
cos[35119]=-78;
cos[35120]=-78;
cos[35121]=-78;
cos[35122]=-78;
cos[35123]=-78;
cos[35124]=-78;
cos[35125]=-78;
cos[35126]=-78;
cos[35127]=-78;
cos[35128]=-78;
cos[35129]=-78;
cos[35130]=-78;
cos[35131]=-78;
cos[35132]=-78;
cos[35133]=-78;
cos[35134]=-78;
cos[35135]=-78;
cos[35136]=-78;
cos[35137]=-78;
cos[35138]=-78;
cos[35139]=-78;
cos[35140]=-78;
cos[35141]=-78;
cos[35142]=-78;
cos[35143]=-78;
cos[35144]=-78;
cos[35145]=-78;
cos[35146]=-78;
cos[35147]=-78;
cos[35148]=-78;
cos[35149]=-78;
cos[35150]=-78;
cos[35151]=-78;
cos[35152]=-78;
cos[35153]=-78;
cos[35154]=-78;
cos[35155]=-78;
cos[35156]=-78;
cos[35157]=-78;
cos[35158]=-78;
cos[35159]=-78;
cos[35160]=-78;
cos[35161]=-78;
cos[35162]=-78;
cos[35163]=-78;
cos[35164]=-78;
cos[35165]=-78;
cos[35166]=-78;
cos[35167]=-78;
cos[35168]=-78;
cos[35169]=-78;
cos[35170]=-78;
cos[35171]=-78;
cos[35172]=-78;
cos[35173]=-78;
cos[35174]=-78;
cos[35175]=-78;
cos[35176]=-78;
cos[35177]=-78;
cos[35178]=-78;
cos[35179]=-78;
cos[35180]=-78;
cos[35181]=-78;
cos[35182]=-78;
cos[35183]=-78;
cos[35184]=-78;
cos[35185]=-78;
cos[35186]=-78;
cos[35187]=-78;
cos[35188]=-78;
cos[35189]=-78;
cos[35190]=-78;
cos[35191]=-78;
cos[35192]=-78;
cos[35193]=-78;
cos[35194]=-78;
cos[35195]=-78;
cos[35196]=-78;
cos[35197]=-78;
cos[35198]=-78;
cos[35199]=-78;
cos[35200]=-78;
cos[35201]=-78;
cos[35202]=-77;
cos[35203]=-77;
cos[35204]=-77;
cos[35205]=-77;
cos[35206]=-77;
cos[35207]=-77;
cos[35208]=-77;
cos[35209]=-77;
cos[35210]=-77;
cos[35211]=-77;
cos[35212]=-77;
cos[35213]=-77;
cos[35214]=-77;
cos[35215]=-77;
cos[35216]=-77;
cos[35217]=-77;
cos[35218]=-77;
cos[35219]=-77;
cos[35220]=-77;
cos[35221]=-77;
cos[35222]=-77;
cos[35223]=-77;
cos[35224]=-77;
cos[35225]=-77;
cos[35226]=-77;
cos[35227]=-77;
cos[35228]=-77;
cos[35229]=-77;
cos[35230]=-77;
cos[35231]=-77;
cos[35232]=-77;
cos[35233]=-77;
cos[35234]=-77;
cos[35235]=-77;
cos[35236]=-77;
cos[35237]=-77;
cos[35238]=-77;
cos[35239]=-77;
cos[35240]=-77;
cos[35241]=-77;
cos[35242]=-77;
cos[35243]=-77;
cos[35244]=-77;
cos[35245]=-77;
cos[35246]=-77;
cos[35247]=-77;
cos[35248]=-77;
cos[35249]=-77;
cos[35250]=-77;
cos[35251]=-77;
cos[35252]=-77;
cos[35253]=-77;
cos[35254]=-77;
cos[35255]=-77;
cos[35256]=-77;
cos[35257]=-77;
cos[35258]=-77;
cos[35259]=-77;
cos[35260]=-77;
cos[35261]=-77;
cos[35262]=-77;
cos[35263]=-77;
cos[35264]=-77;
cos[35265]=-77;
cos[35266]=-77;
cos[35267]=-77;
cos[35268]=-77;
cos[35269]=-77;
cos[35270]=-77;
cos[35271]=-77;
cos[35272]=-77;
cos[35273]=-77;
cos[35274]=-77;
cos[35275]=-77;
cos[35276]=-77;
cos[35277]=-77;
cos[35278]=-77;
cos[35279]=-77;
cos[35280]=-77;
cos[35281]=-77;
cos[35282]=-77;
cos[35283]=-77;
cos[35284]=-77;
cos[35285]=-77;
cos[35286]=-77;
cos[35287]=-77;
cos[35288]=-77;
cos[35289]=-77;
cos[35290]=-77;
cos[35291]=-77;
cos[35292]=-77;
cos[35293]=-77;
cos[35294]=-77;
cos[35295]=-77;
cos[35296]=-77;
cos[35297]=-77;
cos[35298]=-77;
cos[35299]=-77;
cos[35300]=-77;
cos[35301]=-77;
cos[35302]=-77;
cos[35303]=-77;
cos[35304]=-77;
cos[35305]=-77;
cos[35306]=-77;
cos[35307]=-77;
cos[35308]=-77;
cos[35309]=-77;
cos[35310]=-77;
cos[35311]=-77;
cos[35312]=-77;
cos[35313]=-77;
cos[35314]=-77;
cos[35315]=-77;
cos[35316]=-77;
cos[35317]=-77;
cos[35318]=-77;
cos[35319]=-77;
cos[35320]=-77;
cos[35321]=-77;
cos[35322]=-77;
cos[35323]=-77;
cos[35324]=-77;
cos[35325]=-77;
cos[35326]=-76;
cos[35327]=-76;
cos[35328]=-76;
cos[35329]=-76;
cos[35330]=-76;
cos[35331]=-76;
cos[35332]=-76;
cos[35333]=-76;
cos[35334]=-76;
cos[35335]=-76;
cos[35336]=-76;
cos[35337]=-76;
cos[35338]=-76;
cos[35339]=-76;
cos[35340]=-76;
cos[35341]=-76;
cos[35342]=-76;
cos[35343]=-76;
cos[35344]=-76;
cos[35345]=-76;
cos[35346]=-76;
cos[35347]=-76;
cos[35348]=-76;
cos[35349]=-76;
cos[35350]=-76;
cos[35351]=-76;
cos[35352]=-76;
cos[35353]=-76;
cos[35354]=-76;
cos[35355]=-76;
cos[35356]=-76;
cos[35357]=-76;
cos[35358]=-76;
cos[35359]=-76;
cos[35360]=-76;
cos[35361]=-76;
cos[35362]=-76;
cos[35363]=-76;
cos[35364]=-76;
cos[35365]=-76;
cos[35366]=-76;
cos[35367]=-76;
cos[35368]=-76;
cos[35369]=-76;
cos[35370]=-76;
cos[35371]=-76;
cos[35372]=-76;
cos[35373]=-76;
cos[35374]=-76;
cos[35375]=-76;
cos[35376]=-76;
cos[35377]=-76;
cos[35378]=-76;
cos[35379]=-76;
cos[35380]=-76;
cos[35381]=-76;
cos[35382]=-76;
cos[35383]=-76;
cos[35384]=-76;
cos[35385]=-76;
cos[35386]=-76;
cos[35387]=-76;
cos[35388]=-76;
cos[35389]=-76;
cos[35390]=-76;
cos[35391]=-76;
cos[35392]=-76;
cos[35393]=-76;
cos[35394]=-76;
cos[35395]=-76;
cos[35396]=-76;
cos[35397]=-76;
cos[35398]=-76;
cos[35399]=-76;
cos[35400]=-76;
cos[35401]=-76;
cos[35402]=-76;
cos[35403]=-76;
cos[35404]=-76;
cos[35405]=-76;
cos[35406]=-76;
cos[35407]=-76;
cos[35408]=-76;
cos[35409]=-76;
cos[35410]=-76;
cos[35411]=-76;
cos[35412]=-76;
cos[35413]=-76;
cos[35414]=-75;
cos[35415]=-75;
cos[35416]=-75;
cos[35417]=-75;
cos[35418]=-75;
cos[35419]=-75;
cos[35420]=-75;
cos[35421]=-75;
cos[35422]=-75;
cos[35423]=-75;
cos[35424]=-75;
cos[35425]=-75;
cos[35426]=-75;
cos[35427]=-75;
cos[35428]=-75;
cos[35429]=-75;
cos[35430]=-75;
cos[35431]=-75;
cos[35432]=-75;
cos[35433]=-75;
cos[35434]=-75;
cos[35435]=-75;
cos[35436]=-75;
cos[35437]=-75;
cos[35438]=-75;
cos[35439]=-75;
cos[35440]=-75;
cos[35441]=-75;
cos[35442]=-75;
cos[35443]=-75;
cos[35444]=-75;
cos[35445]=-75;
cos[35446]=-75;
cos[35447]=-75;
cos[35448]=-75;
cos[35449]=-75;
cos[35450]=-75;
cos[35451]=-75;
cos[35452]=-75;
cos[35453]=-75;
cos[35454]=-75;
cos[35455]=-75;
cos[35456]=-75;
cos[35457]=-75;
cos[35458]=-75;
cos[35459]=-75;
cos[35460]=-75;
cos[35461]=-75;
cos[35462]=-75;
cos[35463]=-75;
cos[35464]=-75;
cos[35465]=-75;
cos[35466]=-75;
cos[35467]=-75;
cos[35468]=-75;
cos[35469]=-75;
cos[35470]=-75;
cos[35471]=-75;
cos[35472]=-75;
cos[35473]=-75;
cos[35474]=-75;
cos[35475]=-75;
cos[35476]=-75;
cos[35477]=-75;
cos[35478]=-75;
cos[35479]=-75;
cos[35480]=-75;
cos[35481]=-75;
cos[35482]=-75;
cos[35483]=-75;
cos[35484]=-75;
cos[35485]=-75;
cos[35486]=-75;
cos[35487]=-74;
cos[35488]=-74;
cos[35489]=-74;
cos[35490]=-74;
cos[35491]=-74;
cos[35492]=-74;
cos[35493]=-74;
cos[35494]=-74;
cos[35495]=-74;
cos[35496]=-74;
cos[35497]=-74;
cos[35498]=-74;
cos[35499]=-74;
cos[35500]=-74;
cos[35501]=-74;
cos[35502]=-74;
cos[35503]=-74;
cos[35504]=-74;
cos[35505]=-74;
cos[35506]=-74;
cos[35507]=-74;
cos[35508]=-74;
cos[35509]=-74;
cos[35510]=-74;
cos[35511]=-74;
cos[35512]=-74;
cos[35513]=-74;
cos[35514]=-74;
cos[35515]=-74;
cos[35516]=-74;
cos[35517]=-74;
cos[35518]=-74;
cos[35519]=-74;
cos[35520]=-74;
cos[35521]=-74;
cos[35522]=-74;
cos[35523]=-74;
cos[35524]=-74;
cos[35525]=-74;
cos[35526]=-74;
cos[35527]=-74;
cos[35528]=-74;
cos[35529]=-74;
cos[35530]=-74;
cos[35531]=-74;
cos[35532]=-74;
cos[35533]=-74;
cos[35534]=-74;
cos[35535]=-74;
cos[35536]=-74;
cos[35537]=-74;
cos[35538]=-74;
cos[35539]=-74;
cos[35540]=-74;
cos[35541]=-74;
cos[35542]=-74;
cos[35543]=-74;
cos[35544]=-74;
cos[35545]=-74;
cos[35546]=-74;
cos[35547]=-74;
cos[35548]=-74;
cos[35549]=-74;
cos[35550]=-74;
cos[35551]=-73;
cos[35552]=-73;
cos[35553]=-73;
cos[35554]=-73;
cos[35555]=-73;
cos[35556]=-73;
cos[35557]=-73;
cos[35558]=-73;
cos[35559]=-73;
cos[35560]=-73;
cos[35561]=-73;
cos[35562]=-73;
cos[35563]=-73;
cos[35564]=-73;
cos[35565]=-73;
cos[35566]=-73;
cos[35567]=-73;
cos[35568]=-73;
cos[35569]=-73;
cos[35570]=-73;
cos[35571]=-73;
cos[35572]=-73;
cos[35573]=-73;
cos[35574]=-73;
cos[35575]=-73;
cos[35576]=-73;
cos[35577]=-73;
cos[35578]=-73;
cos[35579]=-73;
cos[35580]=-73;
cos[35581]=-73;
cos[35582]=-73;
cos[35583]=-73;
cos[35584]=-73;
cos[35585]=-73;
cos[35586]=-73;
cos[35587]=-73;
cos[35588]=-73;
cos[35589]=-73;
cos[35590]=-73;
cos[35591]=-73;
cos[35592]=-73;
cos[35593]=-73;
cos[35594]=-73;
cos[35595]=-73;
cos[35596]=-73;
cos[35597]=-73;
cos[35598]=-73;
cos[35599]=-73;
cos[35600]=-73;
cos[35601]=-73;
cos[35602]=-73;
cos[35603]=-73;
cos[35604]=-73;
cos[35605]=-73;
cos[35606]=-73;
cos[35607]=-73;
cos[35608]=-72;
cos[35609]=-72;
cos[35610]=-72;
cos[35611]=-72;
cos[35612]=-72;
cos[35613]=-72;
cos[35614]=-72;
cos[35615]=-72;
cos[35616]=-72;
cos[35617]=-72;
cos[35618]=-72;
cos[35619]=-72;
cos[35620]=-72;
cos[35621]=-72;
cos[35622]=-72;
cos[35623]=-72;
cos[35624]=-72;
cos[35625]=-72;
cos[35626]=-72;
cos[35627]=-72;
cos[35628]=-72;
cos[35629]=-72;
cos[35630]=-72;
cos[35631]=-72;
cos[35632]=-72;
cos[35633]=-72;
cos[35634]=-72;
cos[35635]=-72;
cos[35636]=-72;
cos[35637]=-72;
cos[35638]=-72;
cos[35639]=-72;
cos[35640]=-72;
cos[35641]=-72;
cos[35642]=-72;
cos[35643]=-72;
cos[35644]=-72;
cos[35645]=-72;
cos[35646]=-72;
cos[35647]=-72;
cos[35648]=-72;
cos[35649]=-72;
cos[35650]=-72;
cos[35651]=-72;
cos[35652]=-72;
cos[35653]=-72;
cos[35654]=-72;
cos[35655]=-72;
cos[35656]=-72;
cos[35657]=-72;
cos[35658]=-72;
cos[35659]=-72;
cos[35660]=-72;
cos[35661]=-71;
cos[35662]=-71;
cos[35663]=-71;
cos[35664]=-71;
cos[35665]=-71;
cos[35666]=-71;
cos[35667]=-71;
cos[35668]=-71;
cos[35669]=-71;
cos[35670]=-71;
cos[35671]=-71;
cos[35672]=-71;
cos[35673]=-71;
cos[35674]=-71;
cos[35675]=-71;
cos[35676]=-71;
cos[35677]=-71;
cos[35678]=-71;
cos[35679]=-71;
cos[35680]=-71;
cos[35681]=-71;
cos[35682]=-71;
cos[35683]=-71;
cos[35684]=-71;
cos[35685]=-71;
cos[35686]=-71;
cos[35687]=-71;
cos[35688]=-71;
cos[35689]=-71;
cos[35690]=-71;
cos[35691]=-71;
cos[35692]=-71;
cos[35693]=-71;
cos[35694]=-71;
cos[35695]=-71;
cos[35696]=-71;
cos[35697]=-71;
cos[35698]=-71;
cos[35699]=-71;
cos[35700]=-71;
cos[35701]=-71;
cos[35702]=-71;
cos[35703]=-71;
cos[35704]=-71;
cos[35705]=-71;
cos[35706]=-71;
cos[35707]=-71;
cos[35708]=-71;
cos[35709]=-71;
cos[35710]=-70;
cos[35711]=-70;
cos[35712]=-70;
cos[35713]=-70;
cos[35714]=-70;
cos[35715]=-70;
cos[35716]=-70;
cos[35717]=-70;
cos[35718]=-70;
cos[35719]=-70;
cos[35720]=-70;
cos[35721]=-70;
cos[35722]=-70;
cos[35723]=-70;
cos[35724]=-70;
cos[35725]=-70;
cos[35726]=-70;
cos[35727]=-70;
cos[35728]=-70;
cos[35729]=-70;
cos[35730]=-70;
cos[35731]=-70;
cos[35732]=-70;
cos[35733]=-70;
cos[35734]=-70;
cos[35735]=-70;
cos[35736]=-70;
cos[35737]=-70;
cos[35738]=-70;
cos[35739]=-70;
cos[35740]=-70;
cos[35741]=-70;
cos[35742]=-70;
cos[35743]=-70;
cos[35744]=-70;
cos[35745]=-70;
cos[35746]=-70;
cos[35747]=-70;
cos[35748]=-70;
cos[35749]=-70;
cos[35750]=-70;
cos[35751]=-70;
cos[35752]=-70;
cos[35753]=-70;
cos[35754]=-70;
cos[35755]=-69;
cos[35756]=-69;
cos[35757]=-69;
cos[35758]=-69;
cos[35759]=-69;
cos[35760]=-69;
cos[35761]=-69;
cos[35762]=-69;
cos[35763]=-69;
cos[35764]=-69;
cos[35765]=-69;
cos[35766]=-69;
cos[35767]=-69;
cos[35768]=-69;
cos[35769]=-69;
cos[35770]=-69;
cos[35771]=-69;
cos[35772]=-69;
cos[35773]=-69;
cos[35774]=-69;
cos[35775]=-69;
cos[35776]=-69;
cos[35777]=-69;
cos[35778]=-69;
cos[35779]=-69;
cos[35780]=-69;
cos[35781]=-69;
cos[35782]=-69;
cos[35783]=-69;
cos[35784]=-69;
cos[35785]=-69;
cos[35786]=-69;
cos[35787]=-69;
cos[35788]=-69;
cos[35789]=-69;
cos[35790]=-69;
cos[35791]=-69;
cos[35792]=-69;
cos[35793]=-69;
cos[35794]=-69;
cos[35795]=-69;
cos[35796]=-69;
cos[35797]=-69;
cos[35798]=-69;
cos[35799]=-68;
cos[35800]=-68;
cos[35801]=-68;
cos[35802]=-68;
cos[35803]=-68;
cos[35804]=-68;
cos[35805]=-68;
cos[35806]=-68;
cos[35807]=-68;
cos[35808]=-68;
cos[35809]=-68;
cos[35810]=-68;
cos[35811]=-68;
cos[35812]=-68;
cos[35813]=-68;
cos[35814]=-68;
cos[35815]=-68;
cos[35816]=-68;
cos[35817]=-68;
cos[35818]=-68;
cos[35819]=-68;
cos[35820]=-68;
cos[35821]=-68;
cos[35822]=-68;
cos[35823]=-68;
cos[35824]=-68;
cos[35825]=-68;
cos[35826]=-68;
cos[35827]=-68;
cos[35828]=-68;
cos[35829]=-68;
cos[35830]=-68;
cos[35831]=-68;
cos[35832]=-68;
cos[35833]=-68;
cos[35834]=-68;
cos[35835]=-68;
cos[35836]=-68;
cos[35837]=-68;
cos[35838]=-68;
cos[35839]=-68;
cos[35840]=-67;
cos[35841]=-67;
cos[35842]=-67;
cos[35843]=-67;
cos[35844]=-67;
cos[35845]=-67;
cos[35846]=-67;
cos[35847]=-67;
cos[35848]=-67;
cos[35849]=-67;
cos[35850]=-67;
cos[35851]=-67;
cos[35852]=-67;
cos[35853]=-67;
cos[35854]=-67;
cos[35855]=-67;
cos[35856]=-67;
cos[35857]=-67;
cos[35858]=-67;
cos[35859]=-67;
cos[35860]=-67;
cos[35861]=-67;
cos[35862]=-67;
cos[35863]=-67;
cos[35864]=-67;
cos[35865]=-67;
cos[35866]=-67;
cos[35867]=-67;
cos[35868]=-67;
cos[35869]=-67;
cos[35870]=-67;
cos[35871]=-67;
cos[35872]=-67;
cos[35873]=-67;
cos[35874]=-67;
cos[35875]=-67;
cos[35876]=-67;
cos[35877]=-67;
cos[35878]=-67;
cos[35879]=-67;
cos[35880]=-66;
cos[35881]=-66;
cos[35882]=-66;
cos[35883]=-66;
cos[35884]=-66;
cos[35885]=-66;
cos[35886]=-66;
cos[35887]=-66;
cos[35888]=-66;
cos[35889]=-66;
cos[35890]=-66;
cos[35891]=-66;
cos[35892]=-66;
cos[35893]=-66;
cos[35894]=-66;
cos[35895]=-66;
cos[35896]=-66;
cos[35897]=-66;
cos[35898]=-66;
cos[35899]=-66;
cos[35900]=-66;
cos[35901]=-66;
cos[35902]=-66;
cos[35903]=-66;
cos[35904]=-66;
cos[35905]=-66;
cos[35906]=-66;
cos[35907]=-66;
cos[35908]=-66;
cos[35909]=-66;
cos[35910]=-66;
cos[35911]=-66;
cos[35912]=-66;
cos[35913]=-66;
cos[35914]=-66;
cos[35915]=-66;
cos[35916]=-66;
cos[35917]=-66;
cos[35918]=-65;
cos[35919]=-65;
cos[35920]=-65;
cos[35921]=-65;
cos[35922]=-65;
cos[35923]=-65;
cos[35924]=-65;
cos[35925]=-65;
cos[35926]=-65;
cos[35927]=-65;
cos[35928]=-65;
cos[35929]=-65;
cos[35930]=-65;
cos[35931]=-65;
cos[35932]=-65;
cos[35933]=-65;
cos[35934]=-65;
cos[35935]=-65;
cos[35936]=-65;
cos[35937]=-65;
cos[35938]=-65;
cos[35939]=-65;
cos[35940]=-65;
cos[35941]=-65;
cos[35942]=-65;
cos[35943]=-65;
cos[35944]=-65;
cos[35945]=-65;
cos[35946]=-65;
cos[35947]=-65;
cos[35948]=-65;
cos[35949]=-65;
cos[35950]=-65;
cos[35951]=-65;
cos[35952]=-65;
cos[35953]=-65;
cos[35954]=-65;
cos[35955]=-64;
cos[35956]=-64;
cos[35957]=-64;
cos[35958]=-64;
cos[35959]=-64;
cos[35960]=-64;
cos[35961]=-64;
cos[35962]=-64;
cos[35963]=-64;
cos[35964]=-64;
cos[35965]=-64;
cos[35966]=-64;
cos[35967]=-64;
cos[35968]=-64;
cos[35969]=-64;
cos[35970]=-64;
cos[35971]=-64;
cos[35972]=-64;
cos[35973]=-64;
cos[35974]=-64;
cos[35975]=-64;
cos[35976]=-64;
cos[35977]=-64;
cos[35978]=-64;
cos[35979]=-64;
cos[35980]=-64;
cos[35981]=-64;
cos[35982]=-64;
cos[35983]=-64;
cos[35984]=-64;
cos[35985]=-64;
cos[35986]=-64;
cos[35987]=-64;
cos[35988]=-64;
cos[35989]=-64;
cos[35990]=-63;
cos[35991]=-63;
cos[35992]=-63;
cos[35993]=-63;
cos[35994]=-63;
cos[35995]=-63;
cos[35996]=-63;
cos[35997]=-63;
cos[35998]=-63;
cos[35999]=-63;
cos[36000]=-63;
cos[36001]=-63;
cos[36002]=-63;
cos[36003]=-63;
cos[36004]=-63;
cos[36005]=-63;
cos[36006]=-63;
cos[36007]=-63;
cos[36008]=-63;
cos[36009]=-63;
cos[36010]=-63;
cos[36011]=-63;
cos[36012]=-63;
cos[36013]=-63;
cos[36014]=-63;
cos[36015]=-63;
cos[36016]=-63;
cos[36017]=-63;
cos[36018]=-63;
cos[36019]=-63;
cos[36020]=-63;
cos[36021]=-63;
cos[36022]=-63;
cos[36023]=-63;
cos[36024]=-63;
cos[36025]=-62;
cos[36026]=-62;
cos[36027]=-62;
cos[36028]=-62;
cos[36029]=-62;
cos[36030]=-62;
cos[36031]=-62;
cos[36032]=-62;
cos[36033]=-62;
cos[36034]=-62;
cos[36035]=-62;
cos[36036]=-62;
cos[36037]=-62;
cos[36038]=-62;
cos[36039]=-62;
cos[36040]=-62;
cos[36041]=-62;
cos[36042]=-62;
cos[36043]=-62;
cos[36044]=-62;
cos[36045]=-62;
cos[36046]=-62;
cos[36047]=-62;
cos[36048]=-62;
cos[36049]=-62;
cos[36050]=-62;
cos[36051]=-62;
cos[36052]=-62;
cos[36053]=-62;
cos[36054]=-62;
cos[36055]=-62;
cos[36056]=-62;
cos[36057]=-62;
cos[36058]=-61;
cos[36059]=-61;
cos[36060]=-61;
cos[36061]=-61;
cos[36062]=-61;
cos[36063]=-61;
cos[36064]=-61;
cos[36065]=-61;
cos[36066]=-61;
cos[36067]=-61;
cos[36068]=-61;
cos[36069]=-61;
cos[36070]=-61;
cos[36071]=-61;
cos[36072]=-61;
cos[36073]=-61;
cos[36074]=-61;
cos[36075]=-61;
cos[36076]=-61;
cos[36077]=-61;
cos[36078]=-61;
cos[36079]=-61;
cos[36080]=-61;
cos[36081]=-61;
cos[36082]=-61;
cos[36083]=-61;
cos[36084]=-61;
cos[36085]=-61;
cos[36086]=-61;
cos[36087]=-61;
cos[36088]=-61;
cos[36089]=-61;
cos[36090]=-61;
cos[36091]=-60;
cos[36092]=-60;
cos[36093]=-60;
cos[36094]=-60;
cos[36095]=-60;
cos[36096]=-60;
cos[36097]=-60;
cos[36098]=-60;
cos[36099]=-60;
cos[36100]=-60;
cos[36101]=-60;
cos[36102]=-60;
cos[36103]=-60;
cos[36104]=-60;
cos[36105]=-60;
cos[36106]=-60;
cos[36107]=-60;
cos[36108]=-60;
cos[36109]=-60;
cos[36110]=-60;
cos[36111]=-60;
cos[36112]=-60;
cos[36113]=-60;
cos[36114]=-60;
cos[36115]=-60;
cos[36116]=-60;
cos[36117]=-60;
cos[36118]=-60;
cos[36119]=-60;
cos[36120]=-60;
cos[36121]=-60;
cos[36122]=-60;
cos[36123]=-59;
cos[36124]=-59;
cos[36125]=-59;
cos[36126]=-59;
cos[36127]=-59;
cos[36128]=-59;
cos[36129]=-59;
cos[36130]=-59;
cos[36131]=-59;
cos[36132]=-59;
cos[36133]=-59;
cos[36134]=-59;
cos[36135]=-59;
cos[36136]=-59;
cos[36137]=-59;
cos[36138]=-59;
cos[36139]=-59;
cos[36140]=-59;
cos[36141]=-59;
cos[36142]=-59;
cos[36143]=-59;
cos[36144]=-59;
cos[36145]=-59;
cos[36146]=-59;
cos[36147]=-59;
cos[36148]=-59;
cos[36149]=-59;
cos[36150]=-59;
cos[36151]=-59;
cos[36152]=-59;
cos[36153]=-59;
cos[36154]=-58;
cos[36155]=-58;
cos[36156]=-58;
cos[36157]=-58;
cos[36158]=-58;
cos[36159]=-58;
cos[36160]=-58;
cos[36161]=-58;
cos[36162]=-58;
cos[36163]=-58;
cos[36164]=-58;
cos[36165]=-58;
cos[36166]=-58;
cos[36167]=-58;
cos[36168]=-58;
cos[36169]=-58;
cos[36170]=-58;
cos[36171]=-58;
cos[36172]=-58;
cos[36173]=-58;
cos[36174]=-58;
cos[36175]=-58;
cos[36176]=-58;
cos[36177]=-58;
cos[36178]=-58;
cos[36179]=-58;
cos[36180]=-58;
cos[36181]=-58;
cos[36182]=-58;
cos[36183]=-58;
cos[36184]=-57;
cos[36185]=-57;
cos[36186]=-57;
cos[36187]=-57;
cos[36188]=-57;
cos[36189]=-57;
cos[36190]=-57;
cos[36191]=-57;
cos[36192]=-57;
cos[36193]=-57;
cos[36194]=-57;
cos[36195]=-57;
cos[36196]=-57;
cos[36197]=-57;
cos[36198]=-57;
cos[36199]=-57;
cos[36200]=-57;
cos[36201]=-57;
cos[36202]=-57;
cos[36203]=-57;
cos[36204]=-57;
cos[36205]=-57;
cos[36206]=-57;
cos[36207]=-57;
cos[36208]=-57;
cos[36209]=-57;
cos[36210]=-57;
cos[36211]=-57;
cos[36212]=-57;
cos[36213]=-57;
cos[36214]=-56;
cos[36215]=-56;
cos[36216]=-56;
cos[36217]=-56;
cos[36218]=-56;
cos[36219]=-56;
cos[36220]=-56;
cos[36221]=-56;
cos[36222]=-56;
cos[36223]=-56;
cos[36224]=-56;
cos[36225]=-56;
cos[36226]=-56;
cos[36227]=-56;
cos[36228]=-56;
cos[36229]=-56;
cos[36230]=-56;
cos[36231]=-56;
cos[36232]=-56;
cos[36233]=-56;
cos[36234]=-56;
cos[36235]=-56;
cos[36236]=-56;
cos[36237]=-56;
cos[36238]=-56;
cos[36239]=-56;
cos[36240]=-56;
cos[36241]=-56;
cos[36242]=-56;
cos[36243]=-55;
cos[36244]=-55;
cos[36245]=-55;
cos[36246]=-55;
cos[36247]=-55;
cos[36248]=-55;
cos[36249]=-55;
cos[36250]=-55;
cos[36251]=-55;
cos[36252]=-55;
cos[36253]=-55;
cos[36254]=-55;
cos[36255]=-55;
cos[36256]=-55;
cos[36257]=-55;
cos[36258]=-55;
cos[36259]=-55;
cos[36260]=-55;
cos[36261]=-55;
cos[36262]=-55;
cos[36263]=-55;
cos[36264]=-55;
cos[36265]=-55;
cos[36266]=-55;
cos[36267]=-55;
cos[36268]=-55;
cos[36269]=-55;
cos[36270]=-55;
cos[36271]=-55;
cos[36272]=-54;
cos[36273]=-54;
cos[36274]=-54;
cos[36275]=-54;
cos[36276]=-54;
cos[36277]=-54;
cos[36278]=-54;
cos[36279]=-54;
cos[36280]=-54;
cos[36281]=-54;
cos[36282]=-54;
cos[36283]=-54;
cos[36284]=-54;
cos[36285]=-54;
cos[36286]=-54;
cos[36287]=-54;
cos[36288]=-54;
cos[36289]=-54;
cos[36290]=-54;
cos[36291]=-54;
cos[36292]=-54;
cos[36293]=-54;
cos[36294]=-54;
cos[36295]=-54;
cos[36296]=-54;
cos[36297]=-54;
cos[36298]=-54;
cos[36299]=-54;
cos[36300]=-53;
cos[36301]=-53;
cos[36302]=-53;
cos[36303]=-53;
cos[36304]=-53;
cos[36305]=-53;
cos[36306]=-53;
cos[36307]=-53;
cos[36308]=-53;
cos[36309]=-53;
cos[36310]=-53;
cos[36311]=-53;
cos[36312]=-53;
cos[36313]=-53;
cos[36314]=-53;
cos[36315]=-53;
cos[36316]=-53;
cos[36317]=-53;
cos[36318]=-53;
cos[36319]=-53;
cos[36320]=-53;
cos[36321]=-53;
cos[36322]=-53;
cos[36323]=-53;
cos[36324]=-53;
cos[36325]=-53;
cos[36326]=-53;
cos[36327]=-53;
cos[36328]=-52;
cos[36329]=-52;
cos[36330]=-52;
cos[36331]=-52;
cos[36332]=-52;
cos[36333]=-52;
cos[36334]=-52;
cos[36335]=-52;
cos[36336]=-52;
cos[36337]=-52;
cos[36338]=-52;
cos[36339]=-52;
cos[36340]=-52;
cos[36341]=-52;
cos[36342]=-52;
cos[36343]=-52;
cos[36344]=-52;
cos[36345]=-52;
cos[36346]=-52;
cos[36347]=-52;
cos[36348]=-52;
cos[36349]=-52;
cos[36350]=-52;
cos[36351]=-52;
cos[36352]=-52;
cos[36353]=-52;
cos[36354]=-52;
cos[36355]=-51;
cos[36356]=-51;
cos[36357]=-51;
cos[36358]=-51;
cos[36359]=-51;
cos[36360]=-51;
cos[36361]=-51;
cos[36362]=-51;
cos[36363]=-51;
cos[36364]=-51;
cos[36365]=-51;
cos[36366]=-51;
cos[36367]=-51;
cos[36368]=-51;
cos[36369]=-51;
cos[36370]=-51;
cos[36371]=-51;
cos[36372]=-51;
cos[36373]=-51;
cos[36374]=-51;
cos[36375]=-51;
cos[36376]=-51;
cos[36377]=-51;
cos[36378]=-51;
cos[36379]=-51;
cos[36380]=-51;
cos[36381]=-51;
cos[36382]=-50;
cos[36383]=-50;
cos[36384]=-50;
cos[36385]=-50;
cos[36386]=-50;
cos[36387]=-50;
cos[36388]=-50;
cos[36389]=-50;
cos[36390]=-50;
cos[36391]=-50;
cos[36392]=-50;
cos[36393]=-50;
cos[36394]=-50;
cos[36395]=-50;
cos[36396]=-50;
cos[36397]=-50;
cos[36398]=-50;
cos[36399]=-50;
cos[36400]=-50;
cos[36401]=-50;
cos[36402]=-50;
cos[36403]=-50;
cos[36404]=-50;
cos[36405]=-50;
cos[36406]=-50;
cos[36407]=-50;
cos[36408]=-49;
cos[36409]=-49;
cos[36410]=-49;
cos[36411]=-49;
cos[36412]=-49;
cos[36413]=-49;
cos[36414]=-49;
cos[36415]=-49;
cos[36416]=-49;
cos[36417]=-49;
cos[36418]=-49;
cos[36419]=-49;
cos[36420]=-49;
cos[36421]=-49;
cos[36422]=-49;
cos[36423]=-49;
cos[36424]=-49;
cos[36425]=-49;
cos[36426]=-49;
cos[36427]=-49;
cos[36428]=-49;
cos[36429]=-49;
cos[36430]=-49;
cos[36431]=-49;
cos[36432]=-49;
cos[36433]=-49;
cos[36434]=-49;
cos[36435]=-48;
cos[36436]=-48;
cos[36437]=-48;
cos[36438]=-48;
cos[36439]=-48;
cos[36440]=-48;
cos[36441]=-48;
cos[36442]=-48;
cos[36443]=-48;
cos[36444]=-48;
cos[36445]=-48;
cos[36446]=-48;
cos[36447]=-48;
cos[36448]=-48;
cos[36449]=-48;
cos[36450]=-48;
cos[36451]=-48;
cos[36452]=-48;
cos[36453]=-48;
cos[36454]=-48;
cos[36455]=-48;
cos[36456]=-48;
cos[36457]=-48;
cos[36458]=-48;
cos[36459]=-48;
cos[36460]=-47;
cos[36461]=-47;
cos[36462]=-47;
cos[36463]=-47;
cos[36464]=-47;
cos[36465]=-47;
cos[36466]=-47;
cos[36467]=-47;
cos[36468]=-47;
cos[36469]=-47;
cos[36470]=-47;
cos[36471]=-47;
cos[36472]=-47;
cos[36473]=-47;
cos[36474]=-47;
cos[36475]=-47;
cos[36476]=-47;
cos[36477]=-47;
cos[36478]=-47;
cos[36479]=-47;
cos[36480]=-47;
cos[36481]=-47;
cos[36482]=-47;
cos[36483]=-47;
cos[36484]=-47;
cos[36485]=-47;
cos[36486]=-46;
cos[36487]=-46;
cos[36488]=-46;
cos[36489]=-46;
cos[36490]=-46;
cos[36491]=-46;
cos[36492]=-46;
cos[36493]=-46;
cos[36494]=-46;
cos[36495]=-46;
cos[36496]=-46;
cos[36497]=-46;
cos[36498]=-46;
cos[36499]=-46;
cos[36500]=-46;
cos[36501]=-46;
cos[36502]=-46;
cos[36503]=-46;
cos[36504]=-46;
cos[36505]=-46;
cos[36506]=-46;
cos[36507]=-46;
cos[36508]=-46;
cos[36509]=-46;
cos[36510]=-46;
cos[36511]=-45;
cos[36512]=-45;
cos[36513]=-45;
cos[36514]=-45;
cos[36515]=-45;
cos[36516]=-45;
cos[36517]=-45;
cos[36518]=-45;
cos[36519]=-45;
cos[36520]=-45;
cos[36521]=-45;
cos[36522]=-45;
cos[36523]=-45;
cos[36524]=-45;
cos[36525]=-45;
cos[36526]=-45;
cos[36527]=-45;
cos[36528]=-45;
cos[36529]=-45;
cos[36530]=-45;
cos[36531]=-45;
cos[36532]=-45;
cos[36533]=-45;
cos[36534]=-45;
cos[36535]=-45;
cos[36536]=-44;
cos[36537]=-44;
cos[36538]=-44;
cos[36539]=-44;
cos[36540]=-44;
cos[36541]=-44;
cos[36542]=-44;
cos[36543]=-44;
cos[36544]=-44;
cos[36545]=-44;
cos[36546]=-44;
cos[36547]=-44;
cos[36548]=-44;
cos[36549]=-44;
cos[36550]=-44;
cos[36551]=-44;
cos[36552]=-44;
cos[36553]=-44;
cos[36554]=-44;
cos[36555]=-44;
cos[36556]=-44;
cos[36557]=-44;
cos[36558]=-44;
cos[36559]=-44;
cos[36560]=-44;
cos[36561]=-43;
cos[36562]=-43;
cos[36563]=-43;
cos[36564]=-43;
cos[36565]=-43;
cos[36566]=-43;
cos[36567]=-43;
cos[36568]=-43;
cos[36569]=-43;
cos[36570]=-43;
cos[36571]=-43;
cos[36572]=-43;
cos[36573]=-43;
cos[36574]=-43;
cos[36575]=-43;
cos[36576]=-43;
cos[36577]=-43;
cos[36578]=-43;
cos[36579]=-43;
cos[36580]=-43;
cos[36581]=-43;
cos[36582]=-43;
cos[36583]=-43;
cos[36584]=-43;
cos[36585]=-42;
cos[36586]=-42;
cos[36587]=-42;
cos[36588]=-42;
cos[36589]=-42;
cos[36590]=-42;
cos[36591]=-42;
cos[36592]=-42;
cos[36593]=-42;
cos[36594]=-42;
cos[36595]=-42;
cos[36596]=-42;
cos[36597]=-42;
cos[36598]=-42;
cos[36599]=-42;
cos[36600]=-42;
cos[36601]=-42;
cos[36602]=-42;
cos[36603]=-42;
cos[36604]=-42;
cos[36605]=-42;
cos[36606]=-42;
cos[36607]=-42;
cos[36608]=-42;
cos[36609]=-41;
cos[36610]=-41;
cos[36611]=-41;
cos[36612]=-41;
cos[36613]=-41;
cos[36614]=-41;
cos[36615]=-41;
cos[36616]=-41;
cos[36617]=-41;
cos[36618]=-41;
cos[36619]=-41;
cos[36620]=-41;
cos[36621]=-41;
cos[36622]=-41;
cos[36623]=-41;
cos[36624]=-41;
cos[36625]=-41;
cos[36626]=-41;
cos[36627]=-41;
cos[36628]=-41;
cos[36629]=-41;
cos[36630]=-41;
cos[36631]=-41;
cos[36632]=-41;
cos[36633]=-40;
cos[36634]=-40;
cos[36635]=-40;
cos[36636]=-40;
cos[36637]=-40;
cos[36638]=-40;
cos[36639]=-40;
cos[36640]=-40;
cos[36641]=-40;
cos[36642]=-40;
cos[36643]=-40;
cos[36644]=-40;
cos[36645]=-40;
cos[36646]=-40;
cos[36647]=-40;
cos[36648]=-40;
cos[36649]=-40;
cos[36650]=-40;
cos[36651]=-40;
cos[36652]=-40;
cos[36653]=-40;
cos[36654]=-40;
cos[36655]=-40;
cos[36656]=-40;
cos[36657]=-39;
cos[36658]=-39;
cos[36659]=-39;
cos[36660]=-39;
cos[36661]=-39;
cos[36662]=-39;
cos[36663]=-39;
cos[36664]=-39;
cos[36665]=-39;
cos[36666]=-39;
cos[36667]=-39;
cos[36668]=-39;
cos[36669]=-39;
cos[36670]=-39;
cos[36671]=-39;
cos[36672]=-39;
cos[36673]=-39;
cos[36674]=-39;
cos[36675]=-39;
cos[36676]=-39;
cos[36677]=-39;
cos[36678]=-39;
cos[36679]=-39;
cos[36680]=-38;
cos[36681]=-38;
cos[36682]=-38;
cos[36683]=-38;
cos[36684]=-38;
cos[36685]=-38;
cos[36686]=-38;
cos[36687]=-38;
cos[36688]=-38;
cos[36689]=-38;
cos[36690]=-38;
cos[36691]=-38;
cos[36692]=-38;
cos[36693]=-38;
cos[36694]=-38;
cos[36695]=-38;
cos[36696]=-38;
cos[36697]=-38;
cos[36698]=-38;
cos[36699]=-38;
cos[36700]=-38;
cos[36701]=-38;
cos[36702]=-38;
cos[36703]=-38;
cos[36704]=-37;
cos[36705]=-37;
cos[36706]=-37;
cos[36707]=-37;
cos[36708]=-37;
cos[36709]=-37;
cos[36710]=-37;
cos[36711]=-37;
cos[36712]=-37;
cos[36713]=-37;
cos[36714]=-37;
cos[36715]=-37;
cos[36716]=-37;
cos[36717]=-37;
cos[36718]=-37;
cos[36719]=-37;
cos[36720]=-37;
cos[36721]=-37;
cos[36722]=-37;
cos[36723]=-37;
cos[36724]=-37;
cos[36725]=-37;
cos[36726]=-37;
cos[36727]=-36;
cos[36728]=-36;
cos[36729]=-36;
cos[36730]=-36;
cos[36731]=-36;
cos[36732]=-36;
cos[36733]=-36;
cos[36734]=-36;
cos[36735]=-36;
cos[36736]=-36;
cos[36737]=-36;
cos[36738]=-36;
cos[36739]=-36;
cos[36740]=-36;
cos[36741]=-36;
cos[36742]=-36;
cos[36743]=-36;
cos[36744]=-36;
cos[36745]=-36;
cos[36746]=-36;
cos[36747]=-36;
cos[36748]=-36;
cos[36749]=-36;
cos[36750]=-35;
cos[36751]=-35;
cos[36752]=-35;
cos[36753]=-35;
cos[36754]=-35;
cos[36755]=-35;
cos[36756]=-35;
cos[36757]=-35;
cos[36758]=-35;
cos[36759]=-35;
cos[36760]=-35;
cos[36761]=-35;
cos[36762]=-35;
cos[36763]=-35;
cos[36764]=-35;
cos[36765]=-35;
cos[36766]=-35;
cos[36767]=-35;
cos[36768]=-35;
cos[36769]=-35;
cos[36770]=-35;
cos[36771]=-35;
cos[36772]=-35;
cos[36773]=-34;
cos[36774]=-34;
cos[36775]=-34;
cos[36776]=-34;
cos[36777]=-34;
cos[36778]=-34;
cos[36779]=-34;
cos[36780]=-34;
cos[36781]=-34;
cos[36782]=-34;
cos[36783]=-34;
cos[36784]=-34;
cos[36785]=-34;
cos[36786]=-34;
cos[36787]=-34;
cos[36788]=-34;
cos[36789]=-34;
cos[36790]=-34;
cos[36791]=-34;
cos[36792]=-34;
cos[36793]=-34;
cos[36794]=-34;
cos[36795]=-33;
cos[36796]=-33;
cos[36797]=-33;
cos[36798]=-33;
cos[36799]=-33;
cos[36800]=-33;
cos[36801]=-33;
cos[36802]=-33;
cos[36803]=-33;
cos[36804]=-33;
cos[36805]=-33;
cos[36806]=-33;
cos[36807]=-33;
cos[36808]=-33;
cos[36809]=-33;
cos[36810]=-33;
cos[36811]=-33;
cos[36812]=-33;
cos[36813]=-33;
cos[36814]=-33;
cos[36815]=-33;
cos[36816]=-33;
cos[36817]=-33;
cos[36818]=-32;
cos[36819]=-32;
cos[36820]=-32;
cos[36821]=-32;
cos[36822]=-32;
cos[36823]=-32;
cos[36824]=-32;
cos[36825]=-32;
cos[36826]=-32;
cos[36827]=-32;
cos[36828]=-32;
cos[36829]=-32;
cos[36830]=-32;
cos[36831]=-32;
cos[36832]=-32;
cos[36833]=-32;
cos[36834]=-32;
cos[36835]=-32;
cos[36836]=-32;
cos[36837]=-32;
cos[36838]=-32;
cos[36839]=-32;
cos[36840]=-31;
cos[36841]=-31;
cos[36842]=-31;
cos[36843]=-31;
cos[36844]=-31;
cos[36845]=-31;
cos[36846]=-31;
cos[36847]=-31;
cos[36848]=-31;
cos[36849]=-31;
cos[36850]=-31;
cos[36851]=-31;
cos[36852]=-31;
cos[36853]=-31;
cos[36854]=-31;
cos[36855]=-31;
cos[36856]=-31;
cos[36857]=-31;
cos[36858]=-31;
cos[36859]=-31;
cos[36860]=-31;
cos[36861]=-31;
cos[36862]=-30;
cos[36863]=-30;
cos[36864]=-30;
cos[36865]=-30;
cos[36866]=-30;
cos[36867]=-30;
cos[36868]=-30;
cos[36869]=-30;
cos[36870]=-30;
cos[36871]=-30;
cos[36872]=-30;
cos[36873]=-30;
cos[36874]=-30;
cos[36875]=-30;
cos[36876]=-30;
cos[36877]=-30;
cos[36878]=-30;
cos[36879]=-30;
cos[36880]=-30;
cos[36881]=-30;
cos[36882]=-30;
cos[36883]=-30;
cos[36884]=-29;
cos[36885]=-29;
cos[36886]=-29;
cos[36887]=-29;
cos[36888]=-29;
cos[36889]=-29;
cos[36890]=-29;
cos[36891]=-29;
cos[36892]=-29;
cos[36893]=-29;
cos[36894]=-29;
cos[36895]=-29;
cos[36896]=-29;
cos[36897]=-29;
cos[36898]=-29;
cos[36899]=-29;
cos[36900]=-29;
cos[36901]=-29;
cos[36902]=-29;
cos[36903]=-29;
cos[36904]=-29;
cos[36905]=-29;
cos[36906]=-28;
cos[36907]=-28;
cos[36908]=-28;
cos[36909]=-28;
cos[36910]=-28;
cos[36911]=-28;
cos[36912]=-28;
cos[36913]=-28;
cos[36914]=-28;
cos[36915]=-28;
cos[36916]=-28;
cos[36917]=-28;
cos[36918]=-28;
cos[36919]=-28;
cos[36920]=-28;
cos[36921]=-28;
cos[36922]=-28;
cos[36923]=-28;
cos[36924]=-28;
cos[36925]=-28;
cos[36926]=-28;
cos[36927]=-28;
cos[36928]=-27;
cos[36929]=-27;
cos[36930]=-27;
cos[36931]=-27;
cos[36932]=-27;
cos[36933]=-27;
cos[36934]=-27;
cos[36935]=-27;
cos[36936]=-27;
cos[36937]=-27;
cos[36938]=-27;
cos[36939]=-27;
cos[36940]=-27;
cos[36941]=-27;
cos[36942]=-27;
cos[36943]=-27;
cos[36944]=-27;
cos[36945]=-27;
cos[36946]=-27;
cos[36947]=-27;
cos[36948]=-27;
cos[36949]=-27;
cos[36950]=-26;
cos[36951]=-26;
cos[36952]=-26;
cos[36953]=-26;
cos[36954]=-26;
cos[36955]=-26;
cos[36956]=-26;
cos[36957]=-26;
cos[36958]=-26;
cos[36959]=-26;
cos[36960]=-26;
cos[36961]=-26;
cos[36962]=-26;
cos[36963]=-26;
cos[36964]=-26;
cos[36965]=-26;
cos[36966]=-26;
cos[36967]=-26;
cos[36968]=-26;
cos[36969]=-26;
cos[36970]=-26;
cos[36971]=-25;
cos[36972]=-25;
cos[36973]=-25;
cos[36974]=-25;
cos[36975]=-25;
cos[36976]=-25;
cos[36977]=-25;
cos[36978]=-25;
cos[36979]=-25;
cos[36980]=-25;
cos[36981]=-25;
cos[36982]=-25;
cos[36983]=-25;
cos[36984]=-25;
cos[36985]=-25;
cos[36986]=-25;
cos[36987]=-25;
cos[36988]=-25;
cos[36989]=-25;
cos[36990]=-25;
cos[36991]=-25;
cos[36992]=-25;
cos[36993]=-24;
cos[36994]=-24;
cos[36995]=-24;
cos[36996]=-24;
cos[36997]=-24;
cos[36998]=-24;
cos[36999]=-24;
cos[37000]=-24;
cos[37001]=-24;
cos[37002]=-24;
cos[37003]=-24;
cos[37004]=-24;
cos[37005]=-24;
cos[37006]=-24;
cos[37007]=-24;
cos[37008]=-24;
cos[37009]=-24;
cos[37010]=-24;
cos[37011]=-24;
cos[37012]=-24;
cos[37013]=-24;
cos[37014]=-23;
cos[37015]=-23;
cos[37016]=-23;
cos[37017]=-23;
cos[37018]=-23;
cos[37019]=-23;
cos[37020]=-23;
cos[37021]=-23;
cos[37022]=-23;
cos[37023]=-23;
cos[37024]=-23;
cos[37025]=-23;
cos[37026]=-23;
cos[37027]=-23;
cos[37028]=-23;
cos[37029]=-23;
cos[37030]=-23;
cos[37031]=-23;
cos[37032]=-23;
cos[37033]=-23;
cos[37034]=-23;
cos[37035]=-23;
cos[37036]=-22;
cos[37037]=-22;
cos[37038]=-22;
cos[37039]=-22;
cos[37040]=-22;
cos[37041]=-22;
cos[37042]=-22;
cos[37043]=-22;
cos[37044]=-22;
cos[37045]=-22;
cos[37046]=-22;
cos[37047]=-22;
cos[37048]=-22;
cos[37049]=-22;
cos[37050]=-22;
cos[37051]=-22;
cos[37052]=-22;
cos[37053]=-22;
cos[37054]=-22;
cos[37055]=-22;
cos[37056]=-22;
cos[37057]=-21;
cos[37058]=-21;
cos[37059]=-21;
cos[37060]=-21;
cos[37061]=-21;
cos[37062]=-21;
cos[37063]=-21;
cos[37064]=-21;
cos[37065]=-21;
cos[37066]=-21;
cos[37067]=-21;
cos[37068]=-21;
cos[37069]=-21;
cos[37070]=-21;
cos[37071]=-21;
cos[37072]=-21;
cos[37073]=-21;
cos[37074]=-21;
cos[37075]=-21;
cos[37076]=-21;
cos[37077]=-21;
cos[37078]=-20;
cos[37079]=-20;
cos[37080]=-20;
cos[37081]=-20;
cos[37082]=-20;
cos[37083]=-20;
cos[37084]=-20;
cos[37085]=-20;
cos[37086]=-20;
cos[37087]=-20;
cos[37088]=-20;
cos[37089]=-20;
cos[37090]=-20;
cos[37091]=-20;
cos[37092]=-20;
cos[37093]=-20;
cos[37094]=-20;
cos[37095]=-20;
cos[37096]=-20;
cos[37097]=-20;
cos[37098]=-20;
cos[37099]=-19;
cos[37100]=-19;
cos[37101]=-19;
cos[37102]=-19;
cos[37103]=-19;
cos[37104]=-19;
cos[37105]=-19;
cos[37106]=-19;
cos[37107]=-19;
cos[37108]=-19;
cos[37109]=-19;
cos[37110]=-19;
cos[37111]=-19;
cos[37112]=-19;
cos[37113]=-19;
cos[37114]=-19;
cos[37115]=-19;
cos[37116]=-19;
cos[37117]=-19;
cos[37118]=-19;
cos[37119]=-19;
cos[37120]=-18;
cos[37121]=-18;
cos[37122]=-18;
cos[37123]=-18;
cos[37124]=-18;
cos[37125]=-18;
cos[37126]=-18;
cos[37127]=-18;
cos[37128]=-18;
cos[37129]=-18;
cos[37130]=-18;
cos[37131]=-18;
cos[37132]=-18;
cos[37133]=-18;
cos[37134]=-18;
cos[37135]=-18;
cos[37136]=-18;
cos[37137]=-18;
cos[37138]=-18;
cos[37139]=-18;
cos[37140]=-18;
cos[37141]=-17;
cos[37142]=-17;
cos[37143]=-17;
cos[37144]=-17;
cos[37145]=-17;
cos[37146]=-17;
cos[37147]=-17;
cos[37148]=-17;
cos[37149]=-17;
cos[37150]=-17;
cos[37151]=-17;
cos[37152]=-17;
cos[37153]=-17;
cos[37154]=-17;
cos[37155]=-17;
cos[37156]=-17;
cos[37157]=-17;
cos[37158]=-17;
cos[37159]=-17;
cos[37160]=-17;
cos[37161]=-17;
cos[37162]=-16;
cos[37163]=-16;
cos[37164]=-16;
cos[37165]=-16;
cos[37166]=-16;
cos[37167]=-16;
cos[37168]=-16;
cos[37169]=-16;
cos[37170]=-16;
cos[37171]=-16;
cos[37172]=-16;
cos[37173]=-16;
cos[37174]=-16;
cos[37175]=-16;
cos[37176]=-16;
cos[37177]=-16;
cos[37178]=-16;
cos[37179]=-16;
cos[37180]=-16;
cos[37181]=-16;
cos[37182]=-16;
cos[37183]=-15;
cos[37184]=-15;
cos[37185]=-15;
cos[37186]=-15;
cos[37187]=-15;
cos[37188]=-15;
cos[37189]=-15;
cos[37190]=-15;
cos[37191]=-15;
cos[37192]=-15;
cos[37193]=-15;
cos[37194]=-15;
cos[37195]=-15;
cos[37196]=-15;
cos[37197]=-15;
cos[37198]=-15;
cos[37199]=-15;
cos[37200]=-15;
cos[37201]=-15;
cos[37202]=-15;
cos[37203]=-14;
cos[37204]=-14;
cos[37205]=-14;
cos[37206]=-14;
cos[37207]=-14;
cos[37208]=-14;
cos[37209]=-14;
cos[37210]=-14;
cos[37211]=-14;
cos[37212]=-14;
cos[37213]=-14;
cos[37214]=-14;
cos[37215]=-14;
cos[37216]=-14;
cos[37217]=-14;
cos[37218]=-14;
cos[37219]=-14;
cos[37220]=-14;
cos[37221]=-14;
cos[37222]=-14;
cos[37223]=-14;
cos[37224]=-13;
cos[37225]=-13;
cos[37226]=-13;
cos[37227]=-13;
cos[37228]=-13;
cos[37229]=-13;
cos[37230]=-13;
cos[37231]=-13;
cos[37232]=-13;
cos[37233]=-13;
cos[37234]=-13;
cos[37235]=-13;
cos[37236]=-13;
cos[37237]=-13;
cos[37238]=-13;
cos[37239]=-13;
cos[37240]=-13;
cos[37241]=-13;
cos[37242]=-13;
cos[37243]=-13;
cos[37244]=-13;
cos[37245]=-12;
cos[37246]=-12;
cos[37247]=-12;
cos[37248]=-12;
cos[37249]=-12;
cos[37250]=-12;
cos[37251]=-12;
cos[37252]=-12;
cos[37253]=-12;
cos[37254]=-12;
cos[37255]=-12;
cos[37256]=-12;
cos[37257]=-12;
cos[37258]=-12;
cos[37259]=-12;
cos[37260]=-12;
cos[37261]=-12;
cos[37262]=-12;
cos[37263]=-12;
cos[37264]=-12;
cos[37265]=-11;
cos[37266]=-11;
cos[37267]=-11;
cos[37268]=-11;
cos[37269]=-11;
cos[37270]=-11;
cos[37271]=-11;
cos[37272]=-11;
cos[37273]=-11;
cos[37274]=-11;
cos[37275]=-11;
cos[37276]=-11;
cos[37277]=-11;
cos[37278]=-11;
cos[37279]=-11;
cos[37280]=-11;
cos[37281]=-11;
cos[37282]=-11;
cos[37283]=-11;
cos[37284]=-11;
cos[37285]=-11;
cos[37286]=-10;
cos[37287]=-10;
cos[37288]=-10;
cos[37289]=-10;
cos[37290]=-10;
cos[37291]=-10;
cos[37292]=-10;
cos[37293]=-10;
cos[37294]=-10;
cos[37295]=-10;
cos[37296]=-10;
cos[37297]=-10;
cos[37298]=-10;
cos[37299]=-10;
cos[37300]=-10;
cos[37301]=-10;
cos[37302]=-10;
cos[37303]=-10;
cos[37304]=-10;
cos[37305]=-10;
cos[37306]=-9;
cos[37307]=-9;
cos[37308]=-9;
cos[37309]=-9;
cos[37310]=-9;
cos[37311]=-9;
cos[37312]=-9;
cos[37313]=-9;
cos[37314]=-9;
cos[37315]=-9;
cos[37316]=-9;
cos[37317]=-9;
cos[37318]=-9;
cos[37319]=-9;
cos[37320]=-9;
cos[37321]=-9;
cos[37322]=-9;
cos[37323]=-9;
cos[37324]=-9;
cos[37325]=-9;
cos[37326]=-9;
cos[37327]=-8;
cos[37328]=-8;
cos[37329]=-8;
cos[37330]=-8;
cos[37331]=-8;
cos[37332]=-8;
cos[37333]=-8;
cos[37334]=-8;
cos[37335]=-8;
cos[37336]=-8;
cos[37337]=-8;
cos[37338]=-8;
cos[37339]=-8;
cos[37340]=-8;
cos[37341]=-8;
cos[37342]=-8;
cos[37343]=-8;
cos[37344]=-8;
cos[37345]=-8;
cos[37346]=-8;
cos[37347]=-7;
cos[37348]=-7;
cos[37349]=-7;
cos[37350]=-7;
cos[37351]=-7;
cos[37352]=-7;
cos[37353]=-7;
cos[37354]=-7;
cos[37355]=-7;
cos[37356]=-7;
cos[37357]=-7;
cos[37358]=-7;
cos[37359]=-7;
cos[37360]=-7;
cos[37361]=-7;
cos[37362]=-7;
cos[37363]=-7;
cos[37364]=-7;
cos[37365]=-7;
cos[37366]=-7;
cos[37367]=-7;
cos[37368]=-6;
cos[37369]=-6;
cos[37370]=-6;
cos[37371]=-6;
cos[37372]=-6;
cos[37373]=-6;
cos[37374]=-6;
cos[37375]=-6;
cos[37376]=-6;
cos[37377]=-6;
cos[37378]=-6;
cos[37379]=-6;
cos[37380]=-6;
cos[37381]=-6;
cos[37382]=-6;
cos[37383]=-6;
cos[37384]=-6;
cos[37385]=-6;
cos[37386]=-6;
cos[37387]=-6;
cos[37388]=-5;
cos[37389]=-5;
cos[37390]=-5;
cos[37391]=-5;
cos[37392]=-5;
cos[37393]=-5;
cos[37394]=-5;
cos[37395]=-5;
cos[37396]=-5;
cos[37397]=-5;
cos[37398]=-5;
cos[37399]=-5;
cos[37400]=-5;
cos[37401]=-5;
cos[37402]=-5;
cos[37403]=-5;
cos[37404]=-5;
cos[37405]=-5;
cos[37406]=-5;
cos[37407]=-5;
cos[37408]=-5;
cos[37409]=-4;
cos[37410]=-4;
cos[37411]=-4;
cos[37412]=-4;
cos[37413]=-4;
cos[37414]=-4;
cos[37415]=-4;
cos[37416]=-4;
cos[37417]=-4;
cos[37418]=-4;
cos[37419]=-4;
cos[37420]=-4;
cos[37421]=-4;
cos[37422]=-4;
cos[37423]=-4;
cos[37424]=-4;
cos[37425]=-4;
cos[37426]=-4;
cos[37427]=-4;
cos[37428]=-4;
cos[37429]=-3;
cos[37430]=-3;
cos[37431]=-3;
cos[37432]=-3;
cos[37433]=-3;
cos[37434]=-3;
cos[37435]=-3;
cos[37436]=-3;
cos[37437]=-3;
cos[37438]=-3;
cos[37439]=-3;
cos[37440]=-3;
cos[37441]=-3;
cos[37442]=-3;
cos[37443]=-3;
cos[37444]=-3;
cos[37445]=-3;
cos[37446]=-3;
cos[37447]=-3;
cos[37448]=-3;
cos[37449]=-3;
cos[37450]=-2;
cos[37451]=-2;
cos[37452]=-2;
cos[37453]=-2;
cos[37454]=-2;
cos[37455]=-2;
cos[37456]=-2;
cos[37457]=-2;
cos[37458]=-2;
cos[37459]=-2;
cos[37460]=-2;
cos[37461]=-2;
cos[37462]=-2;
cos[37463]=-2;
cos[37464]=-2;
cos[37465]=-2;
cos[37466]=-2;
cos[37467]=-2;
cos[37468]=-2;
cos[37469]=-2;
cos[37470]=-1;
cos[37471]=-1;
cos[37472]=-1;
cos[37473]=-1;
cos[37474]=-1;
cos[37475]=-1;
cos[37476]=-1;
cos[37477]=-1;
cos[37478]=-1;
cos[37479]=-1;
cos[37480]=-1;
cos[37481]=-1;
cos[37482]=-1;
cos[37483]=-1;
cos[37484]=-1;
cos[37485]=-1;
cos[37486]=-1;
cos[37487]=-1;
cos[37488]=-1;
cos[37489]=-1;
cos[37490]=0;
cos[37491]=0;
cos[37492]=0;
cos[37493]=0;
cos[37494]=0;
cos[37495]=0;
cos[37496]=0;
cos[37497]=0;
cos[37498]=0;
cos[37499]=0;
cos[37500]=0;
cos[37501]=0;
cos[37502]=0;
cos[37503]=0;
cos[37504]=0;
cos[37505]=0;
cos[37506]=0;
cos[37507]=0;
cos[37508]=0;
cos[37509]=0;
cos[37510]=0;
cos[37511]=1;
cos[37512]=1;
cos[37513]=1;
cos[37514]=1;
cos[37515]=1;
cos[37516]=1;
cos[37517]=1;
cos[37518]=1;
cos[37519]=1;
cos[37520]=1;
cos[37521]=1;
cos[37522]=1;
cos[37523]=1;
cos[37524]=1;
cos[37525]=1;
cos[37526]=1;
cos[37527]=1;
cos[37528]=1;
cos[37529]=1;
cos[37530]=1;
cos[37531]=2;
cos[37532]=2;
cos[37533]=2;
cos[37534]=2;
cos[37535]=2;
cos[37536]=2;
cos[37537]=2;
cos[37538]=2;
cos[37539]=2;
cos[37540]=2;
cos[37541]=2;
cos[37542]=2;
cos[37543]=2;
cos[37544]=2;
cos[37545]=2;
cos[37546]=2;
cos[37547]=2;
cos[37548]=2;
cos[37549]=2;
cos[37550]=2;
cos[37551]=3;
cos[37552]=3;
cos[37553]=3;
cos[37554]=3;
cos[37555]=3;
cos[37556]=3;
cos[37557]=3;
cos[37558]=3;
cos[37559]=3;
cos[37560]=3;
cos[37561]=3;
cos[37562]=3;
cos[37563]=3;
cos[37564]=3;
cos[37565]=3;
cos[37566]=3;
cos[37567]=3;
cos[37568]=3;
cos[37569]=3;
cos[37570]=3;
cos[37571]=3;
cos[37572]=4;
cos[37573]=4;
cos[37574]=4;
cos[37575]=4;
cos[37576]=4;
cos[37577]=4;
cos[37578]=4;
cos[37579]=4;
cos[37580]=4;
cos[37581]=4;
cos[37582]=4;
cos[37583]=4;
cos[37584]=4;
cos[37585]=4;
cos[37586]=4;
cos[37587]=4;
cos[37588]=4;
cos[37589]=4;
cos[37590]=4;
cos[37591]=4;
cos[37592]=5;
cos[37593]=5;
cos[37594]=5;
cos[37595]=5;
cos[37596]=5;
cos[37597]=5;
cos[37598]=5;
cos[37599]=5;
cos[37600]=5;
cos[37601]=5;
cos[37602]=5;
cos[37603]=5;
cos[37604]=5;
cos[37605]=5;
cos[37606]=5;
cos[37607]=5;
cos[37608]=5;
cos[37609]=5;
cos[37610]=5;
cos[37611]=5;
cos[37612]=5;
cos[37613]=6;
cos[37614]=6;
cos[37615]=6;
cos[37616]=6;
cos[37617]=6;
cos[37618]=6;
cos[37619]=6;
cos[37620]=6;
cos[37621]=6;
cos[37622]=6;
cos[37623]=6;
cos[37624]=6;
cos[37625]=6;
cos[37626]=6;
cos[37627]=6;
cos[37628]=6;
cos[37629]=6;
cos[37630]=6;
cos[37631]=6;
cos[37632]=6;
cos[37633]=7;
cos[37634]=7;
cos[37635]=7;
cos[37636]=7;
cos[37637]=7;
cos[37638]=7;
cos[37639]=7;
cos[37640]=7;
cos[37641]=7;
cos[37642]=7;
cos[37643]=7;
cos[37644]=7;
cos[37645]=7;
cos[37646]=7;
cos[37647]=7;
cos[37648]=7;
cos[37649]=7;
cos[37650]=7;
cos[37651]=7;
cos[37652]=7;
cos[37653]=7;
cos[37654]=8;
cos[37655]=8;
cos[37656]=8;
cos[37657]=8;
cos[37658]=8;
cos[37659]=8;
cos[37660]=8;
cos[37661]=8;
cos[37662]=8;
cos[37663]=8;
cos[37664]=8;
cos[37665]=8;
cos[37666]=8;
cos[37667]=8;
cos[37668]=8;
cos[37669]=8;
cos[37670]=8;
cos[37671]=8;
cos[37672]=8;
cos[37673]=8;
cos[37674]=9;
cos[37675]=9;
cos[37676]=9;
cos[37677]=9;
cos[37678]=9;
cos[37679]=9;
cos[37680]=9;
cos[37681]=9;
cos[37682]=9;
cos[37683]=9;
cos[37684]=9;
cos[37685]=9;
cos[37686]=9;
cos[37687]=9;
cos[37688]=9;
cos[37689]=9;
cos[37690]=9;
cos[37691]=9;
cos[37692]=9;
cos[37693]=9;
cos[37694]=9;
cos[37695]=10;
cos[37696]=10;
cos[37697]=10;
cos[37698]=10;
cos[37699]=10;
cos[37700]=10;
cos[37701]=10;
cos[37702]=10;
cos[37703]=10;
cos[37704]=10;
cos[37705]=10;
cos[37706]=10;
cos[37707]=10;
cos[37708]=10;
cos[37709]=10;
cos[37710]=10;
cos[37711]=10;
cos[37712]=10;
cos[37713]=10;
cos[37714]=10;
cos[37715]=11;
cos[37716]=11;
cos[37717]=11;
cos[37718]=11;
cos[37719]=11;
cos[37720]=11;
cos[37721]=11;
cos[37722]=11;
cos[37723]=11;
cos[37724]=11;
cos[37725]=11;
cos[37726]=11;
cos[37727]=11;
cos[37728]=11;
cos[37729]=11;
cos[37730]=11;
cos[37731]=11;
cos[37732]=11;
cos[37733]=11;
cos[37734]=11;
cos[37735]=11;
cos[37736]=12;
cos[37737]=12;
cos[37738]=12;
cos[37739]=12;
cos[37740]=12;
cos[37741]=12;
cos[37742]=12;
cos[37743]=12;
cos[37744]=12;
cos[37745]=12;
cos[37746]=12;
cos[37747]=12;
cos[37748]=12;
cos[37749]=12;
cos[37750]=12;
cos[37751]=12;
cos[37752]=12;
cos[37753]=12;
cos[37754]=12;
cos[37755]=12;
cos[37756]=13;
cos[37757]=13;
cos[37758]=13;
cos[37759]=13;
cos[37760]=13;
cos[37761]=13;
cos[37762]=13;
cos[37763]=13;
cos[37764]=13;
cos[37765]=13;
cos[37766]=13;
cos[37767]=13;
cos[37768]=13;
cos[37769]=13;
cos[37770]=13;
cos[37771]=13;
cos[37772]=13;
cos[37773]=13;
cos[37774]=13;
cos[37775]=13;
cos[37776]=13;
cos[37777]=14;
cos[37778]=14;
cos[37779]=14;
cos[37780]=14;
cos[37781]=14;
cos[37782]=14;
cos[37783]=14;
cos[37784]=14;
cos[37785]=14;
cos[37786]=14;
cos[37787]=14;
cos[37788]=14;
cos[37789]=14;
cos[37790]=14;
cos[37791]=14;
cos[37792]=14;
cos[37793]=14;
cos[37794]=14;
cos[37795]=14;
cos[37796]=14;
cos[37797]=14;
cos[37798]=15;
cos[37799]=15;
cos[37800]=15;
cos[37801]=15;
cos[37802]=15;
cos[37803]=15;
cos[37804]=15;
cos[37805]=15;
cos[37806]=15;
cos[37807]=15;
cos[37808]=15;
cos[37809]=15;
cos[37810]=15;
cos[37811]=15;
cos[37812]=15;
cos[37813]=15;
cos[37814]=15;
cos[37815]=15;
cos[37816]=15;
cos[37817]=15;
cos[37818]=16;
cos[37819]=16;
cos[37820]=16;
cos[37821]=16;
cos[37822]=16;
cos[37823]=16;
cos[37824]=16;
cos[37825]=16;
cos[37826]=16;
cos[37827]=16;
cos[37828]=16;
cos[37829]=16;
cos[37830]=16;
cos[37831]=16;
cos[37832]=16;
cos[37833]=16;
cos[37834]=16;
cos[37835]=16;
cos[37836]=16;
cos[37837]=16;
cos[37838]=16;
cos[37839]=17;
cos[37840]=17;
cos[37841]=17;
cos[37842]=17;
cos[37843]=17;
cos[37844]=17;
cos[37845]=17;
cos[37846]=17;
cos[37847]=17;
cos[37848]=17;
cos[37849]=17;
cos[37850]=17;
cos[37851]=17;
cos[37852]=17;
cos[37853]=17;
cos[37854]=17;
cos[37855]=17;
cos[37856]=17;
cos[37857]=17;
cos[37858]=17;
cos[37859]=17;
cos[37860]=18;
cos[37861]=18;
cos[37862]=18;
cos[37863]=18;
cos[37864]=18;
cos[37865]=18;
cos[37866]=18;
cos[37867]=18;
cos[37868]=18;
cos[37869]=18;
cos[37870]=18;
cos[37871]=18;
cos[37872]=18;
cos[37873]=18;
cos[37874]=18;
cos[37875]=18;
cos[37876]=18;
cos[37877]=18;
cos[37878]=18;
cos[37879]=18;
cos[37880]=18;
cos[37881]=19;
cos[37882]=19;
cos[37883]=19;
cos[37884]=19;
cos[37885]=19;
cos[37886]=19;
cos[37887]=19;
cos[37888]=19;
cos[37889]=19;
cos[37890]=19;
cos[37891]=19;
cos[37892]=19;
cos[37893]=19;
cos[37894]=19;
cos[37895]=19;
cos[37896]=19;
cos[37897]=19;
cos[37898]=19;
cos[37899]=19;
cos[37900]=19;
cos[37901]=19;
cos[37902]=20;
cos[37903]=20;
cos[37904]=20;
cos[37905]=20;
cos[37906]=20;
cos[37907]=20;
cos[37908]=20;
cos[37909]=20;
cos[37910]=20;
cos[37911]=20;
cos[37912]=20;
cos[37913]=20;
cos[37914]=20;
cos[37915]=20;
cos[37916]=20;
cos[37917]=20;
cos[37918]=20;
cos[37919]=20;
cos[37920]=20;
cos[37921]=20;
cos[37922]=20;
cos[37923]=21;
cos[37924]=21;
cos[37925]=21;
cos[37926]=21;
cos[37927]=21;
cos[37928]=21;
cos[37929]=21;
cos[37930]=21;
cos[37931]=21;
cos[37932]=21;
cos[37933]=21;
cos[37934]=21;
cos[37935]=21;
cos[37936]=21;
cos[37937]=21;
cos[37938]=21;
cos[37939]=21;
cos[37940]=21;
cos[37941]=21;
cos[37942]=21;
cos[37943]=21;
cos[37944]=22;
cos[37945]=22;
cos[37946]=22;
cos[37947]=22;
cos[37948]=22;
cos[37949]=22;
cos[37950]=22;
cos[37951]=22;
cos[37952]=22;
cos[37953]=22;
cos[37954]=22;
cos[37955]=22;
cos[37956]=22;
cos[37957]=22;
cos[37958]=22;
cos[37959]=22;
cos[37960]=22;
cos[37961]=22;
cos[37962]=22;
cos[37963]=22;
cos[37964]=22;
cos[37965]=23;
cos[37966]=23;
cos[37967]=23;
cos[37968]=23;
cos[37969]=23;
cos[37970]=23;
cos[37971]=23;
cos[37972]=23;
cos[37973]=23;
cos[37974]=23;
cos[37975]=23;
cos[37976]=23;
cos[37977]=23;
cos[37978]=23;
cos[37979]=23;
cos[37980]=23;
cos[37981]=23;
cos[37982]=23;
cos[37983]=23;
cos[37984]=23;
cos[37985]=23;
cos[37986]=23;
cos[37987]=24;
cos[37988]=24;
cos[37989]=24;
cos[37990]=24;
cos[37991]=24;
cos[37992]=24;
cos[37993]=24;
cos[37994]=24;
cos[37995]=24;
cos[37996]=24;
cos[37997]=24;
cos[37998]=24;
cos[37999]=24;
cos[38000]=24;
cos[38001]=24;
cos[38002]=24;
cos[38003]=24;
cos[38004]=24;
cos[38005]=24;
cos[38006]=24;
cos[38007]=24;
cos[38008]=25;
cos[38009]=25;
cos[38010]=25;
cos[38011]=25;
cos[38012]=25;
cos[38013]=25;
cos[38014]=25;
cos[38015]=25;
cos[38016]=25;
cos[38017]=25;
cos[38018]=25;
cos[38019]=25;
cos[38020]=25;
cos[38021]=25;
cos[38022]=25;
cos[38023]=25;
cos[38024]=25;
cos[38025]=25;
cos[38026]=25;
cos[38027]=25;
cos[38028]=25;
cos[38029]=25;
cos[38030]=26;
cos[38031]=26;
cos[38032]=26;
cos[38033]=26;
cos[38034]=26;
cos[38035]=26;
cos[38036]=26;
cos[38037]=26;
cos[38038]=26;
cos[38039]=26;
cos[38040]=26;
cos[38041]=26;
cos[38042]=26;
cos[38043]=26;
cos[38044]=26;
cos[38045]=26;
cos[38046]=26;
cos[38047]=26;
cos[38048]=26;
cos[38049]=26;
cos[38050]=26;
cos[38051]=27;
cos[38052]=27;
cos[38053]=27;
cos[38054]=27;
cos[38055]=27;
cos[38056]=27;
cos[38057]=27;
cos[38058]=27;
cos[38059]=27;
cos[38060]=27;
cos[38061]=27;
cos[38062]=27;
cos[38063]=27;
cos[38064]=27;
cos[38065]=27;
cos[38066]=27;
cos[38067]=27;
cos[38068]=27;
cos[38069]=27;
cos[38070]=27;
cos[38071]=27;
cos[38072]=27;
cos[38073]=28;
cos[38074]=28;
cos[38075]=28;
cos[38076]=28;
cos[38077]=28;
cos[38078]=28;
cos[38079]=28;
cos[38080]=28;
cos[38081]=28;
cos[38082]=28;
cos[38083]=28;
cos[38084]=28;
cos[38085]=28;
cos[38086]=28;
cos[38087]=28;
cos[38088]=28;
cos[38089]=28;
cos[38090]=28;
cos[38091]=28;
cos[38092]=28;
cos[38093]=28;
cos[38094]=28;
cos[38095]=29;
cos[38096]=29;
cos[38097]=29;
cos[38098]=29;
cos[38099]=29;
cos[38100]=29;
cos[38101]=29;
cos[38102]=29;
cos[38103]=29;
cos[38104]=29;
cos[38105]=29;
cos[38106]=29;
cos[38107]=29;
cos[38108]=29;
cos[38109]=29;
cos[38110]=29;
cos[38111]=29;
cos[38112]=29;
cos[38113]=29;
cos[38114]=29;
cos[38115]=29;
cos[38116]=29;
cos[38117]=30;
cos[38118]=30;
cos[38119]=30;
cos[38120]=30;
cos[38121]=30;
cos[38122]=30;
cos[38123]=30;
cos[38124]=30;
cos[38125]=30;
cos[38126]=30;
cos[38127]=30;
cos[38128]=30;
cos[38129]=30;
cos[38130]=30;
cos[38131]=30;
cos[38132]=30;
cos[38133]=30;
cos[38134]=30;
cos[38135]=30;
cos[38136]=30;
cos[38137]=30;
cos[38138]=30;
cos[38139]=31;
cos[38140]=31;
cos[38141]=31;
cos[38142]=31;
cos[38143]=31;
cos[38144]=31;
cos[38145]=31;
cos[38146]=31;
cos[38147]=31;
cos[38148]=31;
cos[38149]=31;
cos[38150]=31;
cos[38151]=31;
cos[38152]=31;
cos[38153]=31;
cos[38154]=31;
cos[38155]=31;
cos[38156]=31;
cos[38157]=31;
cos[38158]=31;
cos[38159]=31;
cos[38160]=31;
cos[38161]=32;
cos[38162]=32;
cos[38163]=32;
cos[38164]=32;
cos[38165]=32;
cos[38166]=32;
cos[38167]=32;
cos[38168]=32;
cos[38169]=32;
cos[38170]=32;
cos[38171]=32;
cos[38172]=32;
cos[38173]=32;
cos[38174]=32;
cos[38175]=32;
cos[38176]=32;
cos[38177]=32;
cos[38178]=32;
cos[38179]=32;
cos[38180]=32;
cos[38181]=32;
cos[38182]=32;
cos[38183]=33;
cos[38184]=33;
cos[38185]=33;
cos[38186]=33;
cos[38187]=33;
cos[38188]=33;
cos[38189]=33;
cos[38190]=33;
cos[38191]=33;
cos[38192]=33;
cos[38193]=33;
cos[38194]=33;
cos[38195]=33;
cos[38196]=33;
cos[38197]=33;
cos[38198]=33;
cos[38199]=33;
cos[38200]=33;
cos[38201]=33;
cos[38202]=33;
cos[38203]=33;
cos[38204]=33;
cos[38205]=33;
cos[38206]=34;
cos[38207]=34;
cos[38208]=34;
cos[38209]=34;
cos[38210]=34;
cos[38211]=34;
cos[38212]=34;
cos[38213]=34;
cos[38214]=34;
cos[38215]=34;
cos[38216]=34;
cos[38217]=34;
cos[38218]=34;
cos[38219]=34;
cos[38220]=34;
cos[38221]=34;
cos[38222]=34;
cos[38223]=34;
cos[38224]=34;
cos[38225]=34;
cos[38226]=34;
cos[38227]=34;
cos[38228]=35;
cos[38229]=35;
cos[38230]=35;
cos[38231]=35;
cos[38232]=35;
cos[38233]=35;
cos[38234]=35;
cos[38235]=35;
cos[38236]=35;
cos[38237]=35;
cos[38238]=35;
cos[38239]=35;
cos[38240]=35;
cos[38241]=35;
cos[38242]=35;
cos[38243]=35;
cos[38244]=35;
cos[38245]=35;
cos[38246]=35;
cos[38247]=35;
cos[38248]=35;
cos[38249]=35;
cos[38250]=35;
cos[38251]=36;
cos[38252]=36;
cos[38253]=36;
cos[38254]=36;
cos[38255]=36;
cos[38256]=36;
cos[38257]=36;
cos[38258]=36;
cos[38259]=36;
cos[38260]=36;
cos[38261]=36;
cos[38262]=36;
cos[38263]=36;
cos[38264]=36;
cos[38265]=36;
cos[38266]=36;
cos[38267]=36;
cos[38268]=36;
cos[38269]=36;
cos[38270]=36;
cos[38271]=36;
cos[38272]=36;
cos[38273]=36;
cos[38274]=37;
cos[38275]=37;
cos[38276]=37;
cos[38277]=37;
cos[38278]=37;
cos[38279]=37;
cos[38280]=37;
cos[38281]=37;
cos[38282]=37;
cos[38283]=37;
cos[38284]=37;
cos[38285]=37;
cos[38286]=37;
cos[38287]=37;
cos[38288]=37;
cos[38289]=37;
cos[38290]=37;
cos[38291]=37;
cos[38292]=37;
cos[38293]=37;
cos[38294]=37;
cos[38295]=37;
cos[38296]=37;
cos[38297]=38;
cos[38298]=38;
cos[38299]=38;
cos[38300]=38;
cos[38301]=38;
cos[38302]=38;
cos[38303]=38;
cos[38304]=38;
cos[38305]=38;
cos[38306]=38;
cos[38307]=38;
cos[38308]=38;
cos[38309]=38;
cos[38310]=38;
cos[38311]=38;
cos[38312]=38;
cos[38313]=38;
cos[38314]=38;
cos[38315]=38;
cos[38316]=38;
cos[38317]=38;
cos[38318]=38;
cos[38319]=38;
cos[38320]=38;
cos[38321]=39;
cos[38322]=39;
cos[38323]=39;
cos[38324]=39;
cos[38325]=39;
cos[38326]=39;
cos[38327]=39;
cos[38328]=39;
cos[38329]=39;
cos[38330]=39;
cos[38331]=39;
cos[38332]=39;
cos[38333]=39;
cos[38334]=39;
cos[38335]=39;
cos[38336]=39;
cos[38337]=39;
cos[38338]=39;
cos[38339]=39;
cos[38340]=39;
cos[38341]=39;
cos[38342]=39;
cos[38343]=39;
cos[38344]=40;
cos[38345]=40;
cos[38346]=40;
cos[38347]=40;
cos[38348]=40;
cos[38349]=40;
cos[38350]=40;
cos[38351]=40;
cos[38352]=40;
cos[38353]=40;
cos[38354]=40;
cos[38355]=40;
cos[38356]=40;
cos[38357]=40;
cos[38358]=40;
cos[38359]=40;
cos[38360]=40;
cos[38361]=40;
cos[38362]=40;
cos[38363]=40;
cos[38364]=40;
cos[38365]=40;
cos[38366]=40;
cos[38367]=40;
cos[38368]=41;
cos[38369]=41;
cos[38370]=41;
cos[38371]=41;
cos[38372]=41;
cos[38373]=41;
cos[38374]=41;
cos[38375]=41;
cos[38376]=41;
cos[38377]=41;
cos[38378]=41;
cos[38379]=41;
cos[38380]=41;
cos[38381]=41;
cos[38382]=41;
cos[38383]=41;
cos[38384]=41;
cos[38385]=41;
cos[38386]=41;
cos[38387]=41;
cos[38388]=41;
cos[38389]=41;
cos[38390]=41;
cos[38391]=41;
cos[38392]=42;
cos[38393]=42;
cos[38394]=42;
cos[38395]=42;
cos[38396]=42;
cos[38397]=42;
cos[38398]=42;
cos[38399]=42;
cos[38400]=42;
cos[38401]=42;
cos[38402]=42;
cos[38403]=42;
cos[38404]=42;
cos[38405]=42;
cos[38406]=42;
cos[38407]=42;
cos[38408]=42;
cos[38409]=42;
cos[38410]=42;
cos[38411]=42;
cos[38412]=42;
cos[38413]=42;
cos[38414]=42;
cos[38415]=42;
cos[38416]=43;
cos[38417]=43;
cos[38418]=43;
cos[38419]=43;
cos[38420]=43;
cos[38421]=43;
cos[38422]=43;
cos[38423]=43;
cos[38424]=43;
cos[38425]=43;
cos[38426]=43;
cos[38427]=43;
cos[38428]=43;
cos[38429]=43;
cos[38430]=43;
cos[38431]=43;
cos[38432]=43;
cos[38433]=43;
cos[38434]=43;
cos[38435]=43;
cos[38436]=43;
cos[38437]=43;
cos[38438]=43;
cos[38439]=43;
cos[38440]=44;
cos[38441]=44;
cos[38442]=44;
cos[38443]=44;
cos[38444]=44;
cos[38445]=44;
cos[38446]=44;
cos[38447]=44;
cos[38448]=44;
cos[38449]=44;
cos[38450]=44;
cos[38451]=44;
cos[38452]=44;
cos[38453]=44;
cos[38454]=44;
cos[38455]=44;
cos[38456]=44;
cos[38457]=44;
cos[38458]=44;
cos[38459]=44;
cos[38460]=44;
cos[38461]=44;
cos[38462]=44;
cos[38463]=44;
cos[38464]=44;
cos[38465]=45;
cos[38466]=45;
cos[38467]=45;
cos[38468]=45;
cos[38469]=45;
cos[38470]=45;
cos[38471]=45;
cos[38472]=45;
cos[38473]=45;
cos[38474]=45;
cos[38475]=45;
cos[38476]=45;
cos[38477]=45;
cos[38478]=45;
cos[38479]=45;
cos[38480]=45;
cos[38481]=45;
cos[38482]=45;
cos[38483]=45;
cos[38484]=45;
cos[38485]=45;
cos[38486]=45;
cos[38487]=45;
cos[38488]=45;
cos[38489]=45;
cos[38490]=46;
cos[38491]=46;
cos[38492]=46;
cos[38493]=46;
cos[38494]=46;
cos[38495]=46;
cos[38496]=46;
cos[38497]=46;
cos[38498]=46;
cos[38499]=46;
cos[38500]=46;
cos[38501]=46;
cos[38502]=46;
cos[38503]=46;
cos[38504]=46;
cos[38505]=46;
cos[38506]=46;
cos[38507]=46;
cos[38508]=46;
cos[38509]=46;
cos[38510]=46;
cos[38511]=46;
cos[38512]=46;
cos[38513]=46;
cos[38514]=46;
cos[38515]=47;
cos[38516]=47;
cos[38517]=47;
cos[38518]=47;
cos[38519]=47;
cos[38520]=47;
cos[38521]=47;
cos[38522]=47;
cos[38523]=47;
cos[38524]=47;
cos[38525]=47;
cos[38526]=47;
cos[38527]=47;
cos[38528]=47;
cos[38529]=47;
cos[38530]=47;
cos[38531]=47;
cos[38532]=47;
cos[38533]=47;
cos[38534]=47;
cos[38535]=47;
cos[38536]=47;
cos[38537]=47;
cos[38538]=47;
cos[38539]=47;
cos[38540]=47;
cos[38541]=48;
cos[38542]=48;
cos[38543]=48;
cos[38544]=48;
cos[38545]=48;
cos[38546]=48;
cos[38547]=48;
cos[38548]=48;
cos[38549]=48;
cos[38550]=48;
cos[38551]=48;
cos[38552]=48;
cos[38553]=48;
cos[38554]=48;
cos[38555]=48;
cos[38556]=48;
cos[38557]=48;
cos[38558]=48;
cos[38559]=48;
cos[38560]=48;
cos[38561]=48;
cos[38562]=48;
cos[38563]=48;
cos[38564]=48;
cos[38565]=48;
cos[38566]=49;
cos[38567]=49;
cos[38568]=49;
cos[38569]=49;
cos[38570]=49;
cos[38571]=49;
cos[38572]=49;
cos[38573]=49;
cos[38574]=49;
cos[38575]=49;
cos[38576]=49;
cos[38577]=49;
cos[38578]=49;
cos[38579]=49;
cos[38580]=49;
cos[38581]=49;
cos[38582]=49;
cos[38583]=49;
cos[38584]=49;
cos[38585]=49;
cos[38586]=49;
cos[38587]=49;
cos[38588]=49;
cos[38589]=49;
cos[38590]=49;
cos[38591]=49;
cos[38592]=49;
cos[38593]=50;
cos[38594]=50;
cos[38595]=50;
cos[38596]=50;
cos[38597]=50;
cos[38598]=50;
cos[38599]=50;
cos[38600]=50;
cos[38601]=50;
cos[38602]=50;
cos[38603]=50;
cos[38604]=50;
cos[38605]=50;
cos[38606]=50;
cos[38607]=50;
cos[38608]=50;
cos[38609]=50;
cos[38610]=50;
cos[38611]=50;
cos[38612]=50;
cos[38613]=50;
cos[38614]=50;
cos[38615]=50;
cos[38616]=50;
cos[38617]=50;
cos[38618]=50;
cos[38619]=51;
cos[38620]=51;
cos[38621]=51;
cos[38622]=51;
cos[38623]=51;
cos[38624]=51;
cos[38625]=51;
cos[38626]=51;
cos[38627]=51;
cos[38628]=51;
cos[38629]=51;
cos[38630]=51;
cos[38631]=51;
cos[38632]=51;
cos[38633]=51;
cos[38634]=51;
cos[38635]=51;
cos[38636]=51;
cos[38637]=51;
cos[38638]=51;
cos[38639]=51;
cos[38640]=51;
cos[38641]=51;
cos[38642]=51;
cos[38643]=51;
cos[38644]=51;
cos[38645]=51;
cos[38646]=52;
cos[38647]=52;
cos[38648]=52;
cos[38649]=52;
cos[38650]=52;
cos[38651]=52;
cos[38652]=52;
cos[38653]=52;
cos[38654]=52;
cos[38655]=52;
cos[38656]=52;
cos[38657]=52;
cos[38658]=52;
cos[38659]=52;
cos[38660]=52;
cos[38661]=52;
cos[38662]=52;
cos[38663]=52;
cos[38664]=52;
cos[38665]=52;
cos[38666]=52;
cos[38667]=52;
cos[38668]=52;
cos[38669]=52;
cos[38670]=52;
cos[38671]=52;
cos[38672]=52;
cos[38673]=53;
cos[38674]=53;
cos[38675]=53;
cos[38676]=53;
cos[38677]=53;
cos[38678]=53;
cos[38679]=53;
cos[38680]=53;
cos[38681]=53;
cos[38682]=53;
cos[38683]=53;
cos[38684]=53;
cos[38685]=53;
cos[38686]=53;
cos[38687]=53;
cos[38688]=53;
cos[38689]=53;
cos[38690]=53;
cos[38691]=53;
cos[38692]=53;
cos[38693]=53;
cos[38694]=53;
cos[38695]=53;
cos[38696]=53;
cos[38697]=53;
cos[38698]=53;
cos[38699]=53;
cos[38700]=53;
cos[38701]=54;
cos[38702]=54;
cos[38703]=54;
cos[38704]=54;
cos[38705]=54;
cos[38706]=54;
cos[38707]=54;
cos[38708]=54;
cos[38709]=54;
cos[38710]=54;
cos[38711]=54;
cos[38712]=54;
cos[38713]=54;
cos[38714]=54;
cos[38715]=54;
cos[38716]=54;
cos[38717]=54;
cos[38718]=54;
cos[38719]=54;
cos[38720]=54;
cos[38721]=54;
cos[38722]=54;
cos[38723]=54;
cos[38724]=54;
cos[38725]=54;
cos[38726]=54;
cos[38727]=54;
cos[38728]=54;
cos[38729]=55;
cos[38730]=55;
cos[38731]=55;
cos[38732]=55;
cos[38733]=55;
cos[38734]=55;
cos[38735]=55;
cos[38736]=55;
cos[38737]=55;
cos[38738]=55;
cos[38739]=55;
cos[38740]=55;
cos[38741]=55;
cos[38742]=55;
cos[38743]=55;
cos[38744]=55;
cos[38745]=55;
cos[38746]=55;
cos[38747]=55;
cos[38748]=55;
cos[38749]=55;
cos[38750]=55;
cos[38751]=55;
cos[38752]=55;
cos[38753]=55;
cos[38754]=55;
cos[38755]=55;
cos[38756]=55;
cos[38757]=55;
cos[38758]=56;
cos[38759]=56;
cos[38760]=56;
cos[38761]=56;
cos[38762]=56;
cos[38763]=56;
cos[38764]=56;
cos[38765]=56;
cos[38766]=56;
cos[38767]=56;
cos[38768]=56;
cos[38769]=56;
cos[38770]=56;
cos[38771]=56;
cos[38772]=56;
cos[38773]=56;
cos[38774]=56;
cos[38775]=56;
cos[38776]=56;
cos[38777]=56;
cos[38778]=56;
cos[38779]=56;
cos[38780]=56;
cos[38781]=56;
cos[38782]=56;
cos[38783]=56;
cos[38784]=56;
cos[38785]=56;
cos[38786]=56;
cos[38787]=57;
cos[38788]=57;
cos[38789]=57;
cos[38790]=57;
cos[38791]=57;
cos[38792]=57;
cos[38793]=57;
cos[38794]=57;
cos[38795]=57;
cos[38796]=57;
cos[38797]=57;
cos[38798]=57;
cos[38799]=57;
cos[38800]=57;
cos[38801]=57;
cos[38802]=57;
cos[38803]=57;
cos[38804]=57;
cos[38805]=57;
cos[38806]=57;
cos[38807]=57;
cos[38808]=57;
cos[38809]=57;
cos[38810]=57;
cos[38811]=57;
cos[38812]=57;
cos[38813]=57;
cos[38814]=57;
cos[38815]=57;
cos[38816]=57;
cos[38817]=58;
cos[38818]=58;
cos[38819]=58;
cos[38820]=58;
cos[38821]=58;
cos[38822]=58;
cos[38823]=58;
cos[38824]=58;
cos[38825]=58;
cos[38826]=58;
cos[38827]=58;
cos[38828]=58;
cos[38829]=58;
cos[38830]=58;
cos[38831]=58;
cos[38832]=58;
cos[38833]=58;
cos[38834]=58;
cos[38835]=58;
cos[38836]=58;
cos[38837]=58;
cos[38838]=58;
cos[38839]=58;
cos[38840]=58;
cos[38841]=58;
cos[38842]=58;
cos[38843]=58;
cos[38844]=58;
cos[38845]=58;
cos[38846]=58;
cos[38847]=59;
cos[38848]=59;
cos[38849]=59;
cos[38850]=59;
cos[38851]=59;
cos[38852]=59;
cos[38853]=59;
cos[38854]=59;
cos[38855]=59;
cos[38856]=59;
cos[38857]=59;
cos[38858]=59;
cos[38859]=59;
cos[38860]=59;
cos[38861]=59;
cos[38862]=59;
cos[38863]=59;
cos[38864]=59;
cos[38865]=59;
cos[38866]=59;
cos[38867]=59;
cos[38868]=59;
cos[38869]=59;
cos[38870]=59;
cos[38871]=59;
cos[38872]=59;
cos[38873]=59;
cos[38874]=59;
cos[38875]=59;
cos[38876]=59;
cos[38877]=59;
cos[38878]=60;
cos[38879]=60;
cos[38880]=60;
cos[38881]=60;
cos[38882]=60;
cos[38883]=60;
cos[38884]=60;
cos[38885]=60;
cos[38886]=60;
cos[38887]=60;
cos[38888]=60;
cos[38889]=60;
cos[38890]=60;
cos[38891]=60;
cos[38892]=60;
cos[38893]=60;
cos[38894]=60;
cos[38895]=60;
cos[38896]=60;
cos[38897]=60;
cos[38898]=60;
cos[38899]=60;
cos[38900]=60;
cos[38901]=60;
cos[38902]=60;
cos[38903]=60;
cos[38904]=60;
cos[38905]=60;
cos[38906]=60;
cos[38907]=60;
cos[38908]=60;
cos[38909]=60;
cos[38910]=61;
cos[38911]=61;
cos[38912]=61;
cos[38913]=61;
cos[38914]=61;
cos[38915]=61;
cos[38916]=61;
cos[38917]=61;
cos[38918]=61;
cos[38919]=61;
cos[38920]=61;
cos[38921]=61;
cos[38922]=61;
cos[38923]=61;
cos[38924]=61;
cos[38925]=61;
cos[38926]=61;
cos[38927]=61;
cos[38928]=61;
cos[38929]=61;
cos[38930]=61;
cos[38931]=61;
cos[38932]=61;
cos[38933]=61;
cos[38934]=61;
cos[38935]=61;
cos[38936]=61;
cos[38937]=61;
cos[38938]=61;
cos[38939]=61;
cos[38940]=61;
cos[38941]=61;
cos[38942]=61;
cos[38943]=62;
cos[38944]=62;
cos[38945]=62;
cos[38946]=62;
cos[38947]=62;
cos[38948]=62;
cos[38949]=62;
cos[38950]=62;
cos[38951]=62;
cos[38952]=62;
cos[38953]=62;
cos[38954]=62;
cos[38955]=62;
cos[38956]=62;
cos[38957]=62;
cos[38958]=62;
cos[38959]=62;
cos[38960]=62;
cos[38961]=62;
cos[38962]=62;
cos[38963]=62;
cos[38964]=62;
cos[38965]=62;
cos[38966]=62;
cos[38967]=62;
cos[38968]=62;
cos[38969]=62;
cos[38970]=62;
cos[38971]=62;
cos[38972]=62;
cos[38973]=62;
cos[38974]=62;
cos[38975]=62;
cos[38976]=63;
cos[38977]=63;
cos[38978]=63;
cos[38979]=63;
cos[38980]=63;
cos[38981]=63;
cos[38982]=63;
cos[38983]=63;
cos[38984]=63;
cos[38985]=63;
cos[38986]=63;
cos[38987]=63;
cos[38988]=63;
cos[38989]=63;
cos[38990]=63;
cos[38991]=63;
cos[38992]=63;
cos[38993]=63;
cos[38994]=63;
cos[38995]=63;
cos[38996]=63;
cos[38997]=63;
cos[38998]=63;
cos[38999]=63;
cos[39000]=63;
cos[39001]=63;
cos[39002]=63;
cos[39003]=63;
cos[39004]=63;
cos[39005]=63;
cos[39006]=63;
cos[39007]=63;
cos[39008]=63;
cos[39009]=63;
cos[39010]=63;
cos[39011]=64;
cos[39012]=64;
cos[39013]=64;
cos[39014]=64;
cos[39015]=64;
cos[39016]=64;
cos[39017]=64;
cos[39018]=64;
cos[39019]=64;
cos[39020]=64;
cos[39021]=64;
cos[39022]=64;
cos[39023]=64;
cos[39024]=64;
cos[39025]=64;
cos[39026]=64;
cos[39027]=64;
cos[39028]=64;
cos[39029]=64;
cos[39030]=64;
cos[39031]=64;
cos[39032]=64;
cos[39033]=64;
cos[39034]=64;
cos[39035]=64;
cos[39036]=64;
cos[39037]=64;
cos[39038]=64;
cos[39039]=64;
cos[39040]=64;
cos[39041]=64;
cos[39042]=64;
cos[39043]=64;
cos[39044]=64;
cos[39045]=64;
cos[39046]=65;
cos[39047]=65;
cos[39048]=65;
cos[39049]=65;
cos[39050]=65;
cos[39051]=65;
cos[39052]=65;
cos[39053]=65;
cos[39054]=65;
cos[39055]=65;
cos[39056]=65;
cos[39057]=65;
cos[39058]=65;
cos[39059]=65;
cos[39060]=65;
cos[39061]=65;
cos[39062]=65;
cos[39063]=65;
cos[39064]=65;
cos[39065]=65;
cos[39066]=65;
cos[39067]=65;
cos[39068]=65;
cos[39069]=65;
cos[39070]=65;
cos[39071]=65;
cos[39072]=65;
cos[39073]=65;
cos[39074]=65;
cos[39075]=65;
cos[39076]=65;
cos[39077]=65;
cos[39078]=65;
cos[39079]=65;
cos[39080]=65;
cos[39081]=65;
cos[39082]=65;
cos[39083]=66;
cos[39084]=66;
cos[39085]=66;
cos[39086]=66;
cos[39087]=66;
cos[39088]=66;
cos[39089]=66;
cos[39090]=66;
cos[39091]=66;
cos[39092]=66;
cos[39093]=66;
cos[39094]=66;
cos[39095]=66;
cos[39096]=66;
cos[39097]=66;
cos[39098]=66;
cos[39099]=66;
cos[39100]=66;
cos[39101]=66;
cos[39102]=66;
cos[39103]=66;
cos[39104]=66;
cos[39105]=66;
cos[39106]=66;
cos[39107]=66;
cos[39108]=66;
cos[39109]=66;
cos[39110]=66;
cos[39111]=66;
cos[39112]=66;
cos[39113]=66;
cos[39114]=66;
cos[39115]=66;
cos[39116]=66;
cos[39117]=66;
cos[39118]=66;
cos[39119]=66;
cos[39120]=66;
cos[39121]=67;
cos[39122]=67;
cos[39123]=67;
cos[39124]=67;
cos[39125]=67;
cos[39126]=67;
cos[39127]=67;
cos[39128]=67;
cos[39129]=67;
cos[39130]=67;
cos[39131]=67;
cos[39132]=67;
cos[39133]=67;
cos[39134]=67;
cos[39135]=67;
cos[39136]=67;
cos[39137]=67;
cos[39138]=67;
cos[39139]=67;
cos[39140]=67;
cos[39141]=67;
cos[39142]=67;
cos[39143]=67;
cos[39144]=67;
cos[39145]=67;
cos[39146]=67;
cos[39147]=67;
cos[39148]=67;
cos[39149]=67;
cos[39150]=67;
cos[39151]=67;
cos[39152]=67;
cos[39153]=67;
cos[39154]=67;
cos[39155]=67;
cos[39156]=67;
cos[39157]=67;
cos[39158]=67;
cos[39159]=67;
cos[39160]=67;
cos[39161]=68;
cos[39162]=68;
cos[39163]=68;
cos[39164]=68;
cos[39165]=68;
cos[39166]=68;
cos[39167]=68;
cos[39168]=68;
cos[39169]=68;
cos[39170]=68;
cos[39171]=68;
cos[39172]=68;
cos[39173]=68;
cos[39174]=68;
cos[39175]=68;
cos[39176]=68;
cos[39177]=68;
cos[39178]=68;
cos[39179]=68;
cos[39180]=68;
cos[39181]=68;
cos[39182]=68;
cos[39183]=68;
cos[39184]=68;
cos[39185]=68;
cos[39186]=68;
cos[39187]=68;
cos[39188]=68;
cos[39189]=68;
cos[39190]=68;
cos[39191]=68;
cos[39192]=68;
cos[39193]=68;
cos[39194]=68;
cos[39195]=68;
cos[39196]=68;
cos[39197]=68;
cos[39198]=68;
cos[39199]=68;
cos[39200]=68;
cos[39201]=68;
cos[39202]=69;
cos[39203]=69;
cos[39204]=69;
cos[39205]=69;
cos[39206]=69;
cos[39207]=69;
cos[39208]=69;
cos[39209]=69;
cos[39210]=69;
cos[39211]=69;
cos[39212]=69;
cos[39213]=69;
cos[39214]=69;
cos[39215]=69;
cos[39216]=69;
cos[39217]=69;
cos[39218]=69;
cos[39219]=69;
cos[39220]=69;
cos[39221]=69;
cos[39222]=69;
cos[39223]=69;
cos[39224]=69;
cos[39225]=69;
cos[39226]=69;
cos[39227]=69;
cos[39228]=69;
cos[39229]=69;
cos[39230]=69;
cos[39231]=69;
cos[39232]=69;
cos[39233]=69;
cos[39234]=69;
cos[39235]=69;
cos[39236]=69;
cos[39237]=69;
cos[39238]=69;
cos[39239]=69;
cos[39240]=69;
cos[39241]=69;
cos[39242]=69;
cos[39243]=69;
cos[39244]=69;
cos[39245]=69;
cos[39246]=70;
cos[39247]=70;
cos[39248]=70;
cos[39249]=70;
cos[39250]=70;
cos[39251]=70;
cos[39252]=70;
cos[39253]=70;
cos[39254]=70;
cos[39255]=70;
cos[39256]=70;
cos[39257]=70;
cos[39258]=70;
cos[39259]=70;
cos[39260]=70;
cos[39261]=70;
cos[39262]=70;
cos[39263]=70;
cos[39264]=70;
cos[39265]=70;
cos[39266]=70;
cos[39267]=70;
cos[39268]=70;
cos[39269]=70;
cos[39270]=70;
cos[39271]=70;
cos[39272]=70;
cos[39273]=70;
cos[39274]=70;
cos[39275]=70;
cos[39276]=70;
cos[39277]=70;
cos[39278]=70;
cos[39279]=70;
cos[39280]=70;
cos[39281]=70;
cos[39282]=70;
cos[39283]=70;
cos[39284]=70;
cos[39285]=70;
cos[39286]=70;
cos[39287]=70;
cos[39288]=70;
cos[39289]=70;
cos[39290]=70;
cos[39291]=71;
cos[39292]=71;
cos[39293]=71;
cos[39294]=71;
cos[39295]=71;
cos[39296]=71;
cos[39297]=71;
cos[39298]=71;
cos[39299]=71;
cos[39300]=71;
cos[39301]=71;
cos[39302]=71;
cos[39303]=71;
cos[39304]=71;
cos[39305]=71;
cos[39306]=71;
cos[39307]=71;
cos[39308]=71;
cos[39309]=71;
cos[39310]=71;
cos[39311]=71;
cos[39312]=71;
cos[39313]=71;
cos[39314]=71;
cos[39315]=71;
cos[39316]=71;
cos[39317]=71;
cos[39318]=71;
cos[39319]=71;
cos[39320]=71;
cos[39321]=71;
cos[39322]=71;
cos[39323]=71;
cos[39324]=71;
cos[39325]=71;
cos[39326]=71;
cos[39327]=71;
cos[39328]=71;
cos[39329]=71;
cos[39330]=71;
cos[39331]=71;
cos[39332]=71;
cos[39333]=71;
cos[39334]=71;
cos[39335]=71;
cos[39336]=71;
cos[39337]=71;
cos[39338]=71;
cos[39339]=71;
cos[39340]=72;
cos[39341]=72;
cos[39342]=72;
cos[39343]=72;
cos[39344]=72;
cos[39345]=72;
cos[39346]=72;
cos[39347]=72;
cos[39348]=72;
cos[39349]=72;
cos[39350]=72;
cos[39351]=72;
cos[39352]=72;
cos[39353]=72;
cos[39354]=72;
cos[39355]=72;
cos[39356]=72;
cos[39357]=72;
cos[39358]=72;
cos[39359]=72;
cos[39360]=72;
cos[39361]=72;
cos[39362]=72;
cos[39363]=72;
cos[39364]=72;
cos[39365]=72;
cos[39366]=72;
cos[39367]=72;
cos[39368]=72;
cos[39369]=72;
cos[39370]=72;
cos[39371]=72;
cos[39372]=72;
cos[39373]=72;
cos[39374]=72;
cos[39375]=72;
cos[39376]=72;
cos[39377]=72;
cos[39378]=72;
cos[39379]=72;
cos[39380]=72;
cos[39381]=72;
cos[39382]=72;
cos[39383]=72;
cos[39384]=72;
cos[39385]=72;
cos[39386]=72;
cos[39387]=72;
cos[39388]=72;
cos[39389]=72;
cos[39390]=72;
cos[39391]=72;
cos[39392]=72;
cos[39393]=73;
cos[39394]=73;
cos[39395]=73;
cos[39396]=73;
cos[39397]=73;
cos[39398]=73;
cos[39399]=73;
cos[39400]=73;
cos[39401]=73;
cos[39402]=73;
cos[39403]=73;
cos[39404]=73;
cos[39405]=73;
cos[39406]=73;
cos[39407]=73;
cos[39408]=73;
cos[39409]=73;
cos[39410]=73;
cos[39411]=73;
cos[39412]=73;
cos[39413]=73;
cos[39414]=73;
cos[39415]=73;
cos[39416]=73;
cos[39417]=73;
cos[39418]=73;
cos[39419]=73;
cos[39420]=73;
cos[39421]=73;
cos[39422]=73;
cos[39423]=73;
cos[39424]=73;
cos[39425]=73;
cos[39426]=73;
cos[39427]=73;
cos[39428]=73;
cos[39429]=73;
cos[39430]=73;
cos[39431]=73;
cos[39432]=73;
cos[39433]=73;
cos[39434]=73;
cos[39435]=73;
cos[39436]=73;
cos[39437]=73;
cos[39438]=73;
cos[39439]=73;
cos[39440]=73;
cos[39441]=73;
cos[39442]=73;
cos[39443]=73;
cos[39444]=73;
cos[39445]=73;
cos[39446]=73;
cos[39447]=73;
cos[39448]=73;
cos[39449]=73;
cos[39450]=74;
cos[39451]=74;
cos[39452]=74;
cos[39453]=74;
cos[39454]=74;
cos[39455]=74;
cos[39456]=74;
cos[39457]=74;
cos[39458]=74;
cos[39459]=74;
cos[39460]=74;
cos[39461]=74;
cos[39462]=74;
cos[39463]=74;
cos[39464]=74;
cos[39465]=74;
cos[39466]=74;
cos[39467]=74;
cos[39468]=74;
cos[39469]=74;
cos[39470]=74;
cos[39471]=74;
cos[39472]=74;
cos[39473]=74;
cos[39474]=74;
cos[39475]=74;
cos[39476]=74;
cos[39477]=74;
cos[39478]=74;
cos[39479]=74;
cos[39480]=74;
cos[39481]=74;
cos[39482]=74;
cos[39483]=74;
cos[39484]=74;
cos[39485]=74;
cos[39486]=74;
cos[39487]=74;
cos[39488]=74;
cos[39489]=74;
cos[39490]=74;
cos[39491]=74;
cos[39492]=74;
cos[39493]=74;
cos[39494]=74;
cos[39495]=74;
cos[39496]=74;
cos[39497]=74;
cos[39498]=74;
cos[39499]=74;
cos[39500]=74;
cos[39501]=74;
cos[39502]=74;
cos[39503]=74;
cos[39504]=74;
cos[39505]=74;
cos[39506]=74;
cos[39507]=74;
cos[39508]=74;
cos[39509]=74;
cos[39510]=74;
cos[39511]=74;
cos[39512]=74;
cos[39513]=74;
cos[39514]=75;
cos[39515]=75;
cos[39516]=75;
cos[39517]=75;
cos[39518]=75;
cos[39519]=75;
cos[39520]=75;
cos[39521]=75;
cos[39522]=75;
cos[39523]=75;
cos[39524]=75;
cos[39525]=75;
cos[39526]=75;
cos[39527]=75;
cos[39528]=75;
cos[39529]=75;
cos[39530]=75;
cos[39531]=75;
cos[39532]=75;
cos[39533]=75;
cos[39534]=75;
cos[39535]=75;
cos[39536]=75;
cos[39537]=75;
cos[39538]=75;
cos[39539]=75;
cos[39540]=75;
cos[39541]=75;
cos[39542]=75;
cos[39543]=75;
cos[39544]=75;
cos[39545]=75;
cos[39546]=75;
cos[39547]=75;
cos[39548]=75;
cos[39549]=75;
cos[39550]=75;
cos[39551]=75;
cos[39552]=75;
cos[39553]=75;
cos[39554]=75;
cos[39555]=75;
cos[39556]=75;
cos[39557]=75;
cos[39558]=75;
cos[39559]=75;
cos[39560]=75;
cos[39561]=75;
cos[39562]=75;
cos[39563]=75;
cos[39564]=75;
cos[39565]=75;
cos[39566]=75;
cos[39567]=75;
cos[39568]=75;
cos[39569]=75;
cos[39570]=75;
cos[39571]=75;
cos[39572]=75;
cos[39573]=75;
cos[39574]=75;
cos[39575]=75;
cos[39576]=75;
cos[39577]=75;
cos[39578]=75;
cos[39579]=75;
cos[39580]=75;
cos[39581]=75;
cos[39582]=75;
cos[39583]=75;
cos[39584]=75;
cos[39585]=75;
cos[39586]=75;
cos[39587]=76;
cos[39588]=76;
cos[39589]=76;
cos[39590]=76;
cos[39591]=76;
cos[39592]=76;
cos[39593]=76;
cos[39594]=76;
cos[39595]=76;
cos[39596]=76;
cos[39597]=76;
cos[39598]=76;
cos[39599]=76;
cos[39600]=76;
cos[39601]=76;
cos[39602]=76;
cos[39603]=76;
cos[39604]=76;
cos[39605]=76;
cos[39606]=76;
cos[39607]=76;
cos[39608]=76;
cos[39609]=76;
cos[39610]=76;
cos[39611]=76;
cos[39612]=76;
cos[39613]=76;
cos[39614]=76;
cos[39615]=76;
cos[39616]=76;
cos[39617]=76;
cos[39618]=76;
cos[39619]=76;
cos[39620]=76;
cos[39621]=76;
cos[39622]=76;
cos[39623]=76;
cos[39624]=76;
cos[39625]=76;
cos[39626]=76;
cos[39627]=76;
cos[39628]=76;
cos[39629]=76;
cos[39630]=76;
cos[39631]=76;
cos[39632]=76;
cos[39633]=76;
cos[39634]=76;
cos[39635]=76;
cos[39636]=76;
cos[39637]=76;
cos[39638]=76;
cos[39639]=76;
cos[39640]=76;
cos[39641]=76;
cos[39642]=76;
cos[39643]=76;
cos[39644]=76;
cos[39645]=76;
cos[39646]=76;
cos[39647]=76;
cos[39648]=76;
cos[39649]=76;
cos[39650]=76;
cos[39651]=76;
cos[39652]=76;
cos[39653]=76;
cos[39654]=76;
cos[39655]=76;
cos[39656]=76;
cos[39657]=76;
cos[39658]=76;
cos[39659]=76;
cos[39660]=76;
cos[39661]=76;
cos[39662]=76;
cos[39663]=76;
cos[39664]=76;
cos[39665]=76;
cos[39666]=76;
cos[39667]=76;
cos[39668]=76;
cos[39669]=76;
cos[39670]=76;
cos[39671]=76;
cos[39672]=76;
cos[39673]=76;
cos[39674]=76;
cos[39675]=77;
cos[39676]=77;
cos[39677]=77;
cos[39678]=77;
cos[39679]=77;
cos[39680]=77;
cos[39681]=77;
cos[39682]=77;
cos[39683]=77;
cos[39684]=77;
cos[39685]=77;
cos[39686]=77;
cos[39687]=77;
cos[39688]=77;
cos[39689]=77;
cos[39690]=77;
cos[39691]=77;
cos[39692]=77;
cos[39693]=77;
cos[39694]=77;
cos[39695]=77;
cos[39696]=77;
cos[39697]=77;
cos[39698]=77;
cos[39699]=77;
cos[39700]=77;
cos[39701]=77;
cos[39702]=77;
cos[39703]=77;
cos[39704]=77;
cos[39705]=77;
cos[39706]=77;
cos[39707]=77;
cos[39708]=77;
cos[39709]=77;
cos[39710]=77;
cos[39711]=77;
cos[39712]=77;
cos[39713]=77;
cos[39714]=77;
cos[39715]=77;
cos[39716]=77;
cos[39717]=77;
cos[39718]=77;
cos[39719]=77;
cos[39720]=77;
cos[39721]=77;
cos[39722]=77;
cos[39723]=77;
cos[39724]=77;
cos[39725]=77;
cos[39726]=77;
cos[39727]=77;
cos[39728]=77;
cos[39729]=77;
cos[39730]=77;
cos[39731]=77;
cos[39732]=77;
cos[39733]=77;
cos[39734]=77;
cos[39735]=77;
cos[39736]=77;
cos[39737]=77;
cos[39738]=77;
cos[39739]=77;
cos[39740]=77;
cos[39741]=77;
cos[39742]=77;
cos[39743]=77;
cos[39744]=77;
cos[39745]=77;
cos[39746]=77;
cos[39747]=77;
cos[39748]=77;
cos[39749]=77;
cos[39750]=77;
cos[39751]=77;
cos[39752]=77;
cos[39753]=77;
cos[39754]=77;
cos[39755]=77;
cos[39756]=77;
cos[39757]=77;
cos[39758]=77;
cos[39759]=77;
cos[39760]=77;
cos[39761]=77;
cos[39762]=77;
cos[39763]=77;
cos[39764]=77;
cos[39765]=77;
cos[39766]=77;
cos[39767]=77;
cos[39768]=77;
cos[39769]=77;
cos[39770]=77;
cos[39771]=77;
cos[39772]=77;
cos[39773]=77;
cos[39774]=77;
cos[39775]=77;
cos[39776]=77;
cos[39777]=77;
cos[39778]=77;
cos[39779]=77;
cos[39780]=77;
cos[39781]=77;
cos[39782]=77;
cos[39783]=77;
cos[39784]=77;
cos[39785]=77;
cos[39786]=77;
cos[39787]=77;
cos[39788]=77;
cos[39789]=77;
cos[39790]=77;
cos[39791]=77;
cos[39792]=77;
cos[39793]=77;
cos[39794]=77;
cos[39795]=77;
cos[39796]=77;
cos[39797]=77;
cos[39798]=77;
cos[39799]=78;
cos[39800]=78;
cos[39801]=78;
cos[39802]=78;
cos[39803]=78;
cos[39804]=78;
cos[39805]=78;
cos[39806]=78;
cos[39807]=78;
cos[39808]=78;
cos[39809]=78;
cos[39810]=78;
cos[39811]=78;
cos[39812]=78;
cos[39813]=78;
cos[39814]=78;
cos[39815]=78;
cos[39816]=78;
cos[39817]=78;
cos[39818]=78;
cos[39819]=78;
cos[39820]=78;
cos[39821]=78;
cos[39822]=78;
cos[39823]=78;
cos[39824]=78;
cos[39825]=78;
cos[39826]=78;
cos[39827]=78;
cos[39828]=78;
cos[39829]=78;
cos[39830]=78;
cos[39831]=78;
cos[39832]=78;
cos[39833]=78;
cos[39834]=78;
cos[39835]=78;
cos[39836]=78;
cos[39837]=78;
cos[39838]=78;
cos[39839]=78;
cos[39840]=78;
cos[39841]=78;
cos[39842]=78;
cos[39843]=78;
cos[39844]=78;
cos[39845]=78;
cos[39846]=78;
cos[39847]=78;
cos[39848]=78;
cos[39849]=78;
cos[39850]=78;
cos[39851]=78;
cos[39852]=78;
cos[39853]=78;
cos[39854]=78;
cos[39855]=78;
cos[39856]=78;
cos[39857]=78;
cos[39858]=78;
cos[39859]=78;
cos[39860]=78;
cos[39861]=78;
cos[39862]=78;
cos[39863]=78;
cos[39864]=78;
cos[39865]=78;
cos[39866]=78;
cos[39867]=78;
cos[39868]=78;
cos[39869]=78;
cos[39870]=78;
cos[39871]=78;
cos[39872]=78;
cos[39873]=78;
cos[39874]=78;
cos[39875]=78;
cos[39876]=78;
cos[39877]=78;
cos[39878]=78;
cos[39879]=78;
cos[39880]=78;
cos[39881]=78;
cos[39882]=78;
cos[39883]=78;
cos[39884]=78;
cos[39885]=78;
cos[39886]=78;
cos[39887]=78;
cos[39888]=78;
cos[39889]=78;
cos[39890]=78;
cos[39891]=78;
cos[39892]=78;
cos[39893]=78;
cos[39894]=78;
cos[39895]=78;
cos[39896]=78;
cos[39897]=78;
cos[39898]=78;
cos[39899]=78;
cos[39900]=78;
cos[39901]=78;
cos[39902]=78;
cos[39903]=78;
cos[39904]=78;
cos[39905]=78;
cos[39906]=78;
cos[39907]=78;
cos[39908]=78;
cos[39909]=78;
cos[39910]=78;
cos[39911]=78;
cos[39912]=78;
cos[39913]=78;
cos[39914]=78;
cos[39915]=78;
cos[39916]=78;
cos[39917]=78;
cos[39918]=78;
cos[39919]=78;
cos[39920]=78;
cos[39921]=78;
cos[39922]=78;
cos[39923]=78;
cos[39924]=78;
cos[39925]=78;
cos[39926]=78;
cos[39927]=78;
cos[39928]=78;
cos[39929]=78;
cos[39930]=78;
cos[39931]=78;
cos[39932]=78;
cos[39933]=78;
cos[39934]=78;
cos[39935]=78;
cos[39936]=78;
cos[39937]=78;
cos[39938]=78;
cos[39939]=78;
cos[39940]=78;
cos[39941]=78;
cos[39942]=78;
cos[39943]=78;
cos[39944]=78;
cos[39945]=78;
cos[39946]=78;
cos[39947]=78;
cos[39948]=78;
cos[39949]=78;
cos[39950]=78;
cos[39951]=78;
cos[39952]=78;
cos[39953]=78;
cos[39954]=78;
cos[39955]=78;
cos[39956]=78;
cos[39957]=78;
cos[39958]=78;
cos[39959]=78;
cos[39960]=78;
cos[39961]=78;
cos[39962]=78;
cos[39963]=78;
cos[39964]=78;
cos[39965]=78;
cos[39966]=78;
cos[39967]=78;
cos[39968]=78;
cos[39969]=78;
cos[39970]=78;
cos[39971]=78;
cos[39972]=78;
cos[39973]=78;
cos[39974]=78;
cos[39975]=78;
cos[39976]=78;
cos[39977]=78;
cos[39978]=78;
cos[39979]=78;
cos[39980]=78;
cos[39981]=78;
cos[39982]=78;
cos[39983]=78;
cos[39984]=78;
cos[39985]=78;
cos[39986]=78;
cos[39987]=78;
cos[39988]=78;
cos[39989]=78;
cos[39990]=78;
cos[39991]=78;
cos[39992]=78;
cos[39993]=78;
cos[39994]=78;
cos[39995]=78;
cos[39996]=78;
cos[39997]=78;
cos[39998]=78;
cos[39999]=78;
cos[40000]=78;
sine[0]=0;
sine[1]=0;
sine[2]=0;
sine[3]=0;
sine[4]=0;
sine[5]=0;
sine[6]=0;
sine[7]=0;
sine[8]=0;
sine[9]=0;
sine[10]=0;
sine[11]=1;
sine[12]=1;
sine[13]=1;
sine[14]=1;
sine[15]=1;
sine[16]=1;
sine[17]=1;
sine[18]=1;
sine[19]=1;
sine[20]=1;
sine[21]=1;
sine[22]=1;
sine[23]=1;
sine[24]=1;
sine[25]=1;
sine[26]=1;
sine[27]=1;
sine[28]=1;
sine[29]=1;
sine[30]=1;
sine[31]=2;
sine[32]=2;
sine[33]=2;
sine[34]=2;
sine[35]=2;
sine[36]=2;
sine[37]=2;
sine[38]=2;
sine[39]=2;
sine[40]=2;
sine[41]=2;
sine[42]=2;
sine[43]=2;
sine[44]=2;
sine[45]=2;
sine[46]=2;
sine[47]=2;
sine[48]=2;
sine[49]=2;
sine[50]=2;
sine[51]=3;
sine[52]=3;
sine[53]=3;
sine[54]=3;
sine[55]=3;
sine[56]=3;
sine[57]=3;
sine[58]=3;
sine[59]=3;
sine[60]=3;
sine[61]=3;
sine[62]=3;
sine[63]=3;
sine[64]=3;
sine[65]=3;
sine[66]=3;
sine[67]=3;
sine[68]=3;
sine[69]=3;
sine[70]=3;
sine[71]=3;
sine[72]=4;
sine[73]=4;
sine[74]=4;
sine[75]=4;
sine[76]=4;
sine[77]=4;
sine[78]=4;
sine[79]=4;
sine[80]=4;
sine[81]=4;
sine[82]=4;
sine[83]=4;
sine[84]=4;
sine[85]=4;
sine[86]=4;
sine[87]=4;
sine[88]=4;
sine[89]=4;
sine[90]=4;
sine[91]=4;
sine[92]=5;
sine[93]=5;
sine[94]=5;
sine[95]=5;
sine[96]=5;
sine[97]=5;
sine[98]=5;
sine[99]=5;
sine[100]=5;
sine[101]=5;
sine[102]=5;
sine[103]=5;
sine[104]=5;
sine[105]=5;
sine[106]=5;
sine[107]=5;
sine[108]=5;
sine[109]=5;
sine[110]=5;
sine[111]=5;
sine[112]=5;
sine[113]=6;
sine[114]=6;
sine[115]=6;
sine[116]=6;
sine[117]=6;
sine[118]=6;
sine[119]=6;
sine[120]=6;
sine[121]=6;
sine[122]=6;
sine[123]=6;
sine[124]=6;
sine[125]=6;
sine[126]=6;
sine[127]=6;
sine[128]=6;
sine[129]=6;
sine[130]=6;
sine[131]=6;
sine[132]=6;
sine[133]=7;
sine[134]=7;
sine[135]=7;
sine[136]=7;
sine[137]=7;
sine[138]=7;
sine[139]=7;
sine[140]=7;
sine[141]=7;
sine[142]=7;
sine[143]=7;
sine[144]=7;
sine[145]=7;
sine[146]=7;
sine[147]=7;
sine[148]=7;
sine[149]=7;
sine[150]=7;
sine[151]=7;
sine[152]=7;
sine[153]=7;
sine[154]=8;
sine[155]=8;
sine[156]=8;
sine[157]=8;
sine[158]=8;
sine[159]=8;
sine[160]=8;
sine[161]=8;
sine[162]=8;
sine[163]=8;
sine[164]=8;
sine[165]=8;
sine[166]=8;
sine[167]=8;
sine[168]=8;
sine[169]=8;
sine[170]=8;
sine[171]=8;
sine[172]=8;
sine[173]=8;
sine[174]=9;
sine[175]=9;
sine[176]=9;
sine[177]=9;
sine[178]=9;
sine[179]=9;
sine[180]=9;
sine[181]=9;
sine[182]=9;
sine[183]=9;
sine[184]=9;
sine[185]=9;
sine[186]=9;
sine[187]=9;
sine[188]=9;
sine[189]=9;
sine[190]=9;
sine[191]=9;
sine[192]=9;
sine[193]=9;
sine[194]=9;
sine[195]=10;
sine[196]=10;
sine[197]=10;
sine[198]=10;
sine[199]=10;
sine[200]=10;
sine[201]=10;
sine[202]=10;
sine[203]=10;
sine[204]=10;
sine[205]=10;
sine[206]=10;
sine[207]=10;
sine[208]=10;
sine[209]=10;
sine[210]=10;
sine[211]=10;
sine[212]=10;
sine[213]=10;
sine[214]=10;
sine[215]=11;
sine[216]=11;
sine[217]=11;
sine[218]=11;
sine[219]=11;
sine[220]=11;
sine[221]=11;
sine[222]=11;
sine[223]=11;
sine[224]=11;
sine[225]=11;
sine[226]=11;
sine[227]=11;
sine[228]=11;
sine[229]=11;
sine[230]=11;
sine[231]=11;
sine[232]=11;
sine[233]=11;
sine[234]=11;
sine[235]=11;
sine[236]=12;
sine[237]=12;
sine[238]=12;
sine[239]=12;
sine[240]=12;
sine[241]=12;
sine[242]=12;
sine[243]=12;
sine[244]=12;
sine[245]=12;
sine[246]=12;
sine[247]=12;
sine[248]=12;
sine[249]=12;
sine[250]=12;
sine[251]=12;
sine[252]=12;
sine[253]=12;
sine[254]=12;
sine[255]=12;
sine[256]=13;
sine[257]=13;
sine[258]=13;
sine[259]=13;
sine[260]=13;
sine[261]=13;
sine[262]=13;
sine[263]=13;
sine[264]=13;
sine[265]=13;
sine[266]=13;
sine[267]=13;
sine[268]=13;
sine[269]=13;
sine[270]=13;
sine[271]=13;
sine[272]=13;
sine[273]=13;
sine[274]=13;
sine[275]=13;
sine[276]=13;
sine[277]=14;
sine[278]=14;
sine[279]=14;
sine[280]=14;
sine[281]=14;
sine[282]=14;
sine[283]=14;
sine[284]=14;
sine[285]=14;
sine[286]=14;
sine[287]=14;
sine[288]=14;
sine[289]=14;
sine[290]=14;
sine[291]=14;
sine[292]=14;
sine[293]=14;
sine[294]=14;
sine[295]=14;
sine[296]=14;
sine[297]=14;
sine[298]=15;
sine[299]=15;
sine[300]=15;
sine[301]=15;
sine[302]=15;
sine[303]=15;
sine[304]=15;
sine[305]=15;
sine[306]=15;
sine[307]=15;
sine[308]=15;
sine[309]=15;
sine[310]=15;
sine[311]=15;
sine[312]=15;
sine[313]=15;
sine[314]=15;
sine[315]=15;
sine[316]=15;
sine[317]=15;
sine[318]=16;
sine[319]=16;
sine[320]=16;
sine[321]=16;
sine[322]=16;
sine[323]=16;
sine[324]=16;
sine[325]=16;
sine[326]=16;
sine[327]=16;
sine[328]=16;
sine[329]=16;
sine[330]=16;
sine[331]=16;
sine[332]=16;
sine[333]=16;
sine[334]=16;
sine[335]=16;
sine[336]=16;
sine[337]=16;
sine[338]=16;
sine[339]=17;
sine[340]=17;
sine[341]=17;
sine[342]=17;
sine[343]=17;
sine[344]=17;
sine[345]=17;
sine[346]=17;
sine[347]=17;
sine[348]=17;
sine[349]=17;
sine[350]=17;
sine[351]=17;
sine[352]=17;
sine[353]=17;
sine[354]=17;
sine[355]=17;
sine[356]=17;
sine[357]=17;
sine[358]=17;
sine[359]=17;
sine[360]=18;
sine[361]=18;
sine[362]=18;
sine[363]=18;
sine[364]=18;
sine[365]=18;
sine[366]=18;
sine[367]=18;
sine[368]=18;
sine[369]=18;
sine[370]=18;
sine[371]=18;
sine[372]=18;
sine[373]=18;
sine[374]=18;
sine[375]=18;
sine[376]=18;
sine[377]=18;
sine[378]=18;
sine[379]=18;
sine[380]=18;
sine[381]=19;
sine[382]=19;
sine[383]=19;
sine[384]=19;
sine[385]=19;
sine[386]=19;
sine[387]=19;
sine[388]=19;
sine[389]=19;
sine[390]=19;
sine[391]=19;
sine[392]=19;
sine[393]=19;
sine[394]=19;
sine[395]=19;
sine[396]=19;
sine[397]=19;
sine[398]=19;
sine[399]=19;
sine[400]=19;
sine[401]=19;
sine[402]=20;
sine[403]=20;
sine[404]=20;
sine[405]=20;
sine[406]=20;
sine[407]=20;
sine[408]=20;
sine[409]=20;
sine[410]=20;
sine[411]=20;
sine[412]=20;
sine[413]=20;
sine[414]=20;
sine[415]=20;
sine[416]=20;
sine[417]=20;
sine[418]=20;
sine[419]=20;
sine[420]=20;
sine[421]=20;
sine[422]=20;
sine[423]=21;
sine[424]=21;
sine[425]=21;
sine[426]=21;
sine[427]=21;
sine[428]=21;
sine[429]=21;
sine[430]=21;
sine[431]=21;
sine[432]=21;
sine[433]=21;
sine[434]=21;
sine[435]=21;
sine[436]=21;
sine[437]=21;
sine[438]=21;
sine[439]=21;
sine[440]=21;
sine[441]=21;
sine[442]=21;
sine[443]=21;
sine[444]=22;
sine[445]=22;
sine[446]=22;
sine[447]=22;
sine[448]=22;
sine[449]=22;
sine[450]=22;
sine[451]=22;
sine[452]=22;
sine[453]=22;
sine[454]=22;
sine[455]=22;
sine[456]=22;
sine[457]=22;
sine[458]=22;
sine[459]=22;
sine[460]=22;
sine[461]=22;
sine[462]=22;
sine[463]=22;
sine[464]=22;
sine[465]=23;
sine[466]=23;
sine[467]=23;
sine[468]=23;
sine[469]=23;
sine[470]=23;
sine[471]=23;
sine[472]=23;
sine[473]=23;
sine[474]=23;
sine[475]=23;
sine[476]=23;
sine[477]=23;
sine[478]=23;
sine[479]=23;
sine[480]=23;
sine[481]=23;
sine[482]=23;
sine[483]=23;
sine[484]=23;
sine[485]=23;
sine[486]=23;
sine[487]=24;
sine[488]=24;
sine[489]=24;
sine[490]=24;
sine[491]=24;
sine[492]=24;
sine[493]=24;
sine[494]=24;
sine[495]=24;
sine[496]=24;
sine[497]=24;
sine[498]=24;
sine[499]=24;
sine[500]=24;
sine[501]=24;
sine[502]=24;
sine[503]=24;
sine[504]=24;
sine[505]=24;
sine[506]=24;
sine[507]=24;
sine[508]=25;
sine[509]=25;
sine[510]=25;
sine[511]=25;
sine[512]=25;
sine[513]=25;
sine[514]=25;
sine[515]=25;
sine[516]=25;
sine[517]=25;
sine[518]=25;
sine[519]=25;
sine[520]=25;
sine[521]=25;
sine[522]=25;
sine[523]=25;
sine[524]=25;
sine[525]=25;
sine[526]=25;
sine[527]=25;
sine[528]=25;
sine[529]=25;
sine[530]=26;
sine[531]=26;
sine[532]=26;
sine[533]=26;
sine[534]=26;
sine[535]=26;
sine[536]=26;
sine[537]=26;
sine[538]=26;
sine[539]=26;
sine[540]=26;
sine[541]=26;
sine[542]=26;
sine[543]=26;
sine[544]=26;
sine[545]=26;
sine[546]=26;
sine[547]=26;
sine[548]=26;
sine[549]=26;
sine[550]=26;
sine[551]=27;
sine[552]=27;
sine[553]=27;
sine[554]=27;
sine[555]=27;
sine[556]=27;
sine[557]=27;
sine[558]=27;
sine[559]=27;
sine[560]=27;
sine[561]=27;
sine[562]=27;
sine[563]=27;
sine[564]=27;
sine[565]=27;
sine[566]=27;
sine[567]=27;
sine[568]=27;
sine[569]=27;
sine[570]=27;
sine[571]=27;
sine[572]=27;
sine[573]=28;
sine[574]=28;
sine[575]=28;
sine[576]=28;
sine[577]=28;
sine[578]=28;
sine[579]=28;
sine[580]=28;
sine[581]=28;
sine[582]=28;
sine[583]=28;
sine[584]=28;
sine[585]=28;
sine[586]=28;
sine[587]=28;
sine[588]=28;
sine[589]=28;
sine[590]=28;
sine[591]=28;
sine[592]=28;
sine[593]=28;
sine[594]=28;
sine[595]=29;
sine[596]=29;
sine[597]=29;
sine[598]=29;
sine[599]=29;
sine[600]=29;
sine[601]=29;
sine[602]=29;
sine[603]=29;
sine[604]=29;
sine[605]=29;
sine[606]=29;
sine[607]=29;
sine[608]=29;
sine[609]=29;
sine[610]=29;
sine[611]=29;
sine[612]=29;
sine[613]=29;
sine[614]=29;
sine[615]=29;
sine[616]=29;
sine[617]=30;
sine[618]=30;
sine[619]=30;
sine[620]=30;
sine[621]=30;
sine[622]=30;
sine[623]=30;
sine[624]=30;
sine[625]=30;
sine[626]=30;
sine[627]=30;
sine[628]=30;
sine[629]=30;
sine[630]=30;
sine[631]=30;
sine[632]=30;
sine[633]=30;
sine[634]=30;
sine[635]=30;
sine[636]=30;
sine[637]=30;
sine[638]=30;
sine[639]=31;
sine[640]=31;
sine[641]=31;
sine[642]=31;
sine[643]=31;
sine[644]=31;
sine[645]=31;
sine[646]=31;
sine[647]=31;
sine[648]=31;
sine[649]=31;
sine[650]=31;
sine[651]=31;
sine[652]=31;
sine[653]=31;
sine[654]=31;
sine[655]=31;
sine[656]=31;
sine[657]=31;
sine[658]=31;
sine[659]=31;
sine[660]=31;
sine[661]=32;
sine[662]=32;
sine[663]=32;
sine[664]=32;
sine[665]=32;
sine[666]=32;
sine[667]=32;
sine[668]=32;
sine[669]=32;
sine[670]=32;
sine[671]=32;
sine[672]=32;
sine[673]=32;
sine[674]=32;
sine[675]=32;
sine[676]=32;
sine[677]=32;
sine[678]=32;
sine[679]=32;
sine[680]=32;
sine[681]=32;
sine[682]=32;
sine[683]=33;
sine[684]=33;
sine[685]=33;
sine[686]=33;
sine[687]=33;
sine[688]=33;
sine[689]=33;
sine[690]=33;
sine[691]=33;
sine[692]=33;
sine[693]=33;
sine[694]=33;
sine[695]=33;
sine[696]=33;
sine[697]=33;
sine[698]=33;
sine[699]=33;
sine[700]=33;
sine[701]=33;
sine[702]=33;
sine[703]=33;
sine[704]=33;
sine[705]=33;
sine[706]=34;
sine[707]=34;
sine[708]=34;
sine[709]=34;
sine[710]=34;
sine[711]=34;
sine[712]=34;
sine[713]=34;
sine[714]=34;
sine[715]=34;
sine[716]=34;
sine[717]=34;
sine[718]=34;
sine[719]=34;
sine[720]=34;
sine[721]=34;
sine[722]=34;
sine[723]=34;
sine[724]=34;
sine[725]=34;
sine[726]=34;
sine[727]=34;
sine[728]=35;
sine[729]=35;
sine[730]=35;
sine[731]=35;
sine[732]=35;
sine[733]=35;
sine[734]=35;
sine[735]=35;
sine[736]=35;
sine[737]=35;
sine[738]=35;
sine[739]=35;
sine[740]=35;
sine[741]=35;
sine[742]=35;
sine[743]=35;
sine[744]=35;
sine[745]=35;
sine[746]=35;
sine[747]=35;
sine[748]=35;
sine[749]=35;
sine[750]=35;
sine[751]=36;
sine[752]=36;
sine[753]=36;
sine[754]=36;
sine[755]=36;
sine[756]=36;
sine[757]=36;
sine[758]=36;
sine[759]=36;
sine[760]=36;
sine[761]=36;
sine[762]=36;
sine[763]=36;
sine[764]=36;
sine[765]=36;
sine[766]=36;
sine[767]=36;
sine[768]=36;
sine[769]=36;
sine[770]=36;
sine[771]=36;
sine[772]=36;
sine[773]=36;
sine[774]=37;
sine[775]=37;
sine[776]=37;
sine[777]=37;
sine[778]=37;
sine[779]=37;
sine[780]=37;
sine[781]=37;
sine[782]=37;
sine[783]=37;
sine[784]=37;
sine[785]=37;
sine[786]=37;
sine[787]=37;
sine[788]=37;
sine[789]=37;
sine[790]=37;
sine[791]=37;
sine[792]=37;
sine[793]=37;
sine[794]=37;
sine[795]=37;
sine[796]=37;
sine[797]=38;
sine[798]=38;
sine[799]=38;
sine[800]=38;
sine[801]=38;
sine[802]=38;
sine[803]=38;
sine[804]=38;
sine[805]=38;
sine[806]=38;
sine[807]=38;
sine[808]=38;
sine[809]=38;
sine[810]=38;
sine[811]=38;
sine[812]=38;
sine[813]=38;
sine[814]=38;
sine[815]=38;
sine[816]=38;
sine[817]=38;
sine[818]=38;
sine[819]=38;
sine[820]=38;
sine[821]=39;
sine[822]=39;
sine[823]=39;
sine[824]=39;
sine[825]=39;
sine[826]=39;
sine[827]=39;
sine[828]=39;
sine[829]=39;
sine[830]=39;
sine[831]=39;
sine[832]=39;
sine[833]=39;
sine[834]=39;
sine[835]=39;
sine[836]=39;
sine[837]=39;
sine[838]=39;
sine[839]=39;
sine[840]=39;
sine[841]=39;
sine[842]=39;
sine[843]=39;
sine[844]=40;
sine[845]=40;
sine[846]=40;
sine[847]=40;
sine[848]=40;
sine[849]=40;
sine[850]=40;
sine[851]=40;
sine[852]=40;
sine[853]=40;
sine[854]=40;
sine[855]=40;
sine[856]=40;
sine[857]=40;
sine[858]=40;
sine[859]=40;
sine[860]=40;
sine[861]=40;
sine[862]=40;
sine[863]=40;
sine[864]=40;
sine[865]=40;
sine[866]=40;
sine[867]=40;
sine[868]=41;
sine[869]=41;
sine[870]=41;
sine[871]=41;
sine[872]=41;
sine[873]=41;
sine[874]=41;
sine[875]=41;
sine[876]=41;
sine[877]=41;
sine[878]=41;
sine[879]=41;
sine[880]=41;
sine[881]=41;
sine[882]=41;
sine[883]=41;
sine[884]=41;
sine[885]=41;
sine[886]=41;
sine[887]=41;
sine[888]=41;
sine[889]=41;
sine[890]=41;
sine[891]=41;
sine[892]=42;
sine[893]=42;
sine[894]=42;
sine[895]=42;
sine[896]=42;
sine[897]=42;
sine[898]=42;
sine[899]=42;
sine[900]=42;
sine[901]=42;
sine[902]=42;
sine[903]=42;
sine[904]=42;
sine[905]=42;
sine[906]=42;
sine[907]=42;
sine[908]=42;
sine[909]=42;
sine[910]=42;
sine[911]=42;
sine[912]=42;
sine[913]=42;
sine[914]=42;
sine[915]=42;
sine[916]=43;
sine[917]=43;
sine[918]=43;
sine[919]=43;
sine[920]=43;
sine[921]=43;
sine[922]=43;
sine[923]=43;
sine[924]=43;
sine[925]=43;
sine[926]=43;
sine[927]=43;
sine[928]=43;
sine[929]=43;
sine[930]=43;
sine[931]=43;
sine[932]=43;
sine[933]=43;
sine[934]=43;
sine[935]=43;
sine[936]=43;
sine[937]=43;
sine[938]=43;
sine[939]=43;
sine[940]=44;
sine[941]=44;
sine[942]=44;
sine[943]=44;
sine[944]=44;
sine[945]=44;
sine[946]=44;
sine[947]=44;
sine[948]=44;
sine[949]=44;
sine[950]=44;
sine[951]=44;
sine[952]=44;
sine[953]=44;
sine[954]=44;
sine[955]=44;
sine[956]=44;
sine[957]=44;
sine[958]=44;
sine[959]=44;
sine[960]=44;
sine[961]=44;
sine[962]=44;
sine[963]=44;
sine[964]=44;
sine[965]=45;
sine[966]=45;
sine[967]=45;
sine[968]=45;
sine[969]=45;
sine[970]=45;
sine[971]=45;
sine[972]=45;
sine[973]=45;
sine[974]=45;
sine[975]=45;
sine[976]=45;
sine[977]=45;
sine[978]=45;
sine[979]=45;
sine[980]=45;
sine[981]=45;
sine[982]=45;
sine[983]=45;
sine[984]=45;
sine[985]=45;
sine[986]=45;
sine[987]=45;
sine[988]=45;
sine[989]=45;
sine[990]=46;
sine[991]=46;
sine[992]=46;
sine[993]=46;
sine[994]=46;
sine[995]=46;
sine[996]=46;
sine[997]=46;
sine[998]=46;
sine[999]=46;
sine[1000]=46;
sine[1001]=46;
sine[1002]=46;
sine[1003]=46;
sine[1004]=46;
sine[1005]=46;
sine[1006]=46;
sine[1007]=46;
sine[1008]=46;
sine[1009]=46;
sine[1010]=46;
sine[1011]=46;
sine[1012]=46;
sine[1013]=46;
sine[1014]=46;
sine[1015]=47;
sine[1016]=47;
sine[1017]=47;
sine[1018]=47;
sine[1019]=47;
sine[1020]=47;
sine[1021]=47;
sine[1022]=47;
sine[1023]=47;
sine[1024]=47;
sine[1025]=47;
sine[1026]=47;
sine[1027]=47;
sine[1028]=47;
sine[1029]=47;
sine[1030]=47;
sine[1031]=47;
sine[1032]=47;
sine[1033]=47;
sine[1034]=47;
sine[1035]=47;
sine[1036]=47;
sine[1037]=47;
sine[1038]=47;
sine[1039]=47;
sine[1040]=47;
sine[1041]=48;
sine[1042]=48;
sine[1043]=48;
sine[1044]=48;
sine[1045]=48;
sine[1046]=48;
sine[1047]=48;
sine[1048]=48;
sine[1049]=48;
sine[1050]=48;
sine[1051]=48;
sine[1052]=48;
sine[1053]=48;
sine[1054]=48;
sine[1055]=48;
sine[1056]=48;
sine[1057]=48;
sine[1058]=48;
sine[1059]=48;
sine[1060]=48;
sine[1061]=48;
sine[1062]=48;
sine[1063]=48;
sine[1064]=48;
sine[1065]=48;
sine[1066]=49;
sine[1067]=49;
sine[1068]=49;
sine[1069]=49;
sine[1070]=49;
sine[1071]=49;
sine[1072]=49;
sine[1073]=49;
sine[1074]=49;
sine[1075]=49;
sine[1076]=49;
sine[1077]=49;
sine[1078]=49;
sine[1079]=49;
sine[1080]=49;
sine[1081]=49;
sine[1082]=49;
sine[1083]=49;
sine[1084]=49;
sine[1085]=49;
sine[1086]=49;
sine[1087]=49;
sine[1088]=49;
sine[1089]=49;
sine[1090]=49;
sine[1091]=49;
sine[1092]=49;
sine[1093]=50;
sine[1094]=50;
sine[1095]=50;
sine[1096]=50;
sine[1097]=50;
sine[1098]=50;
sine[1099]=50;
sine[1100]=50;
sine[1101]=50;
sine[1102]=50;
sine[1103]=50;
sine[1104]=50;
sine[1105]=50;
sine[1106]=50;
sine[1107]=50;
sine[1108]=50;
sine[1109]=50;
sine[1110]=50;
sine[1111]=50;
sine[1112]=50;
sine[1113]=50;
sine[1114]=50;
sine[1115]=50;
sine[1116]=50;
sine[1117]=50;
sine[1118]=50;
sine[1119]=51;
sine[1120]=51;
sine[1121]=51;
sine[1122]=51;
sine[1123]=51;
sine[1124]=51;
sine[1125]=51;
sine[1126]=51;
sine[1127]=51;
sine[1128]=51;
sine[1129]=51;
sine[1130]=51;
sine[1131]=51;
sine[1132]=51;
sine[1133]=51;
sine[1134]=51;
sine[1135]=51;
sine[1136]=51;
sine[1137]=51;
sine[1138]=51;
sine[1139]=51;
sine[1140]=51;
sine[1141]=51;
sine[1142]=51;
sine[1143]=51;
sine[1144]=51;
sine[1145]=51;
sine[1146]=52;
sine[1147]=52;
sine[1148]=52;
sine[1149]=52;
sine[1150]=52;
sine[1151]=52;
sine[1152]=52;
sine[1153]=52;
sine[1154]=52;
sine[1155]=52;
sine[1156]=52;
sine[1157]=52;
sine[1158]=52;
sine[1159]=52;
sine[1160]=52;
sine[1161]=52;
sine[1162]=52;
sine[1163]=52;
sine[1164]=52;
sine[1165]=52;
sine[1166]=52;
sine[1167]=52;
sine[1168]=52;
sine[1169]=52;
sine[1170]=52;
sine[1171]=52;
sine[1172]=52;
sine[1173]=53;
sine[1174]=53;
sine[1175]=53;
sine[1176]=53;
sine[1177]=53;
sine[1178]=53;
sine[1179]=53;
sine[1180]=53;
sine[1181]=53;
sine[1182]=53;
sine[1183]=53;
sine[1184]=53;
sine[1185]=53;
sine[1186]=53;
sine[1187]=53;
sine[1188]=53;
sine[1189]=53;
sine[1190]=53;
sine[1191]=53;
sine[1192]=53;
sine[1193]=53;
sine[1194]=53;
sine[1195]=53;
sine[1196]=53;
sine[1197]=53;
sine[1198]=53;
sine[1199]=53;
sine[1200]=53;
sine[1201]=54;
sine[1202]=54;
sine[1203]=54;
sine[1204]=54;
sine[1205]=54;
sine[1206]=54;
sine[1207]=54;
sine[1208]=54;
sine[1209]=54;
sine[1210]=54;
sine[1211]=54;
sine[1212]=54;
sine[1213]=54;
sine[1214]=54;
sine[1215]=54;
sine[1216]=54;
sine[1217]=54;
sine[1218]=54;
sine[1219]=54;
sine[1220]=54;
sine[1221]=54;
sine[1222]=54;
sine[1223]=54;
sine[1224]=54;
sine[1225]=54;
sine[1226]=54;
sine[1227]=54;
sine[1228]=54;
sine[1229]=55;
sine[1230]=55;
sine[1231]=55;
sine[1232]=55;
sine[1233]=55;
sine[1234]=55;
sine[1235]=55;
sine[1236]=55;
sine[1237]=55;
sine[1238]=55;
sine[1239]=55;
sine[1240]=55;
sine[1241]=55;
sine[1242]=55;
sine[1243]=55;
sine[1244]=55;
sine[1245]=55;
sine[1246]=55;
sine[1247]=55;
sine[1248]=55;
sine[1249]=55;
sine[1250]=55;
sine[1251]=55;
sine[1252]=55;
sine[1253]=55;
sine[1254]=55;
sine[1255]=55;
sine[1256]=55;
sine[1257]=55;
sine[1258]=56;
sine[1259]=56;
sine[1260]=56;
sine[1261]=56;
sine[1262]=56;
sine[1263]=56;
sine[1264]=56;
sine[1265]=56;
sine[1266]=56;
sine[1267]=56;
sine[1268]=56;
sine[1269]=56;
sine[1270]=56;
sine[1271]=56;
sine[1272]=56;
sine[1273]=56;
sine[1274]=56;
sine[1275]=56;
sine[1276]=56;
sine[1277]=56;
sine[1278]=56;
sine[1279]=56;
sine[1280]=56;
sine[1281]=56;
sine[1282]=56;
sine[1283]=56;
sine[1284]=56;
sine[1285]=56;
sine[1286]=56;
sine[1287]=57;
sine[1288]=57;
sine[1289]=57;
sine[1290]=57;
sine[1291]=57;
sine[1292]=57;
sine[1293]=57;
sine[1294]=57;
sine[1295]=57;
sine[1296]=57;
sine[1297]=57;
sine[1298]=57;
sine[1299]=57;
sine[1300]=57;
sine[1301]=57;
sine[1302]=57;
sine[1303]=57;
sine[1304]=57;
sine[1305]=57;
sine[1306]=57;
sine[1307]=57;
sine[1308]=57;
sine[1309]=57;
sine[1310]=57;
sine[1311]=57;
sine[1312]=57;
sine[1313]=57;
sine[1314]=57;
sine[1315]=57;
sine[1316]=57;
sine[1317]=58;
sine[1318]=58;
sine[1319]=58;
sine[1320]=58;
sine[1321]=58;
sine[1322]=58;
sine[1323]=58;
sine[1324]=58;
sine[1325]=58;
sine[1326]=58;
sine[1327]=58;
sine[1328]=58;
sine[1329]=58;
sine[1330]=58;
sine[1331]=58;
sine[1332]=58;
sine[1333]=58;
sine[1334]=58;
sine[1335]=58;
sine[1336]=58;
sine[1337]=58;
sine[1338]=58;
sine[1339]=58;
sine[1340]=58;
sine[1341]=58;
sine[1342]=58;
sine[1343]=58;
sine[1344]=58;
sine[1345]=58;
sine[1346]=58;
sine[1347]=59;
sine[1348]=59;
sine[1349]=59;
sine[1350]=59;
sine[1351]=59;
sine[1352]=59;
sine[1353]=59;
sine[1354]=59;
sine[1355]=59;
sine[1356]=59;
sine[1357]=59;
sine[1358]=59;
sine[1359]=59;
sine[1360]=59;
sine[1361]=59;
sine[1362]=59;
sine[1363]=59;
sine[1364]=59;
sine[1365]=59;
sine[1366]=59;
sine[1367]=59;
sine[1368]=59;
sine[1369]=59;
sine[1370]=59;
sine[1371]=59;
sine[1372]=59;
sine[1373]=59;
sine[1374]=59;
sine[1375]=59;
sine[1376]=59;
sine[1377]=59;
sine[1378]=60;
sine[1379]=60;
sine[1380]=60;
sine[1381]=60;
sine[1382]=60;
sine[1383]=60;
sine[1384]=60;
sine[1385]=60;
sine[1386]=60;
sine[1387]=60;
sine[1388]=60;
sine[1389]=60;
sine[1390]=60;
sine[1391]=60;
sine[1392]=60;
sine[1393]=60;
sine[1394]=60;
sine[1395]=60;
sine[1396]=60;
sine[1397]=60;
sine[1398]=60;
sine[1399]=60;
sine[1400]=60;
sine[1401]=60;
sine[1402]=60;
sine[1403]=60;
sine[1404]=60;
sine[1405]=60;
sine[1406]=60;
sine[1407]=60;
sine[1408]=60;
sine[1409]=60;
sine[1410]=61;
sine[1411]=61;
sine[1412]=61;
sine[1413]=61;
sine[1414]=61;
sine[1415]=61;
sine[1416]=61;
sine[1417]=61;
sine[1418]=61;
sine[1419]=61;
sine[1420]=61;
sine[1421]=61;
sine[1422]=61;
sine[1423]=61;
sine[1424]=61;
sine[1425]=61;
sine[1426]=61;
sine[1427]=61;
sine[1428]=61;
sine[1429]=61;
sine[1430]=61;
sine[1431]=61;
sine[1432]=61;
sine[1433]=61;
sine[1434]=61;
sine[1435]=61;
sine[1436]=61;
sine[1437]=61;
sine[1438]=61;
sine[1439]=61;
sine[1440]=61;
sine[1441]=61;
sine[1442]=61;
sine[1443]=62;
sine[1444]=62;
sine[1445]=62;
sine[1446]=62;
sine[1447]=62;
sine[1448]=62;
sine[1449]=62;
sine[1450]=62;
sine[1451]=62;
sine[1452]=62;
sine[1453]=62;
sine[1454]=62;
sine[1455]=62;
sine[1456]=62;
sine[1457]=62;
sine[1458]=62;
sine[1459]=62;
sine[1460]=62;
sine[1461]=62;
sine[1462]=62;
sine[1463]=62;
sine[1464]=62;
sine[1465]=62;
sine[1466]=62;
sine[1467]=62;
sine[1468]=62;
sine[1469]=62;
sine[1470]=62;
sine[1471]=62;
sine[1472]=62;
sine[1473]=62;
sine[1474]=62;
sine[1475]=62;
sine[1476]=63;
sine[1477]=63;
sine[1478]=63;
sine[1479]=63;
sine[1480]=63;
sine[1481]=63;
sine[1482]=63;
sine[1483]=63;
sine[1484]=63;
sine[1485]=63;
sine[1486]=63;
sine[1487]=63;
sine[1488]=63;
sine[1489]=63;
sine[1490]=63;
sine[1491]=63;
sine[1492]=63;
sine[1493]=63;
sine[1494]=63;
sine[1495]=63;
sine[1496]=63;
sine[1497]=63;
sine[1498]=63;
sine[1499]=63;
sine[1500]=63;
sine[1501]=63;
sine[1502]=63;
sine[1503]=63;
sine[1504]=63;
sine[1505]=63;
sine[1506]=63;
sine[1507]=63;
sine[1508]=63;
sine[1509]=63;
sine[1510]=63;
sine[1511]=64;
sine[1512]=64;
sine[1513]=64;
sine[1514]=64;
sine[1515]=64;
sine[1516]=64;
sine[1517]=64;
sine[1518]=64;
sine[1519]=64;
sine[1520]=64;
sine[1521]=64;
sine[1522]=64;
sine[1523]=64;
sine[1524]=64;
sine[1525]=64;
sine[1526]=64;
sine[1527]=64;
sine[1528]=64;
sine[1529]=64;
sine[1530]=64;
sine[1531]=64;
sine[1532]=64;
sine[1533]=64;
sine[1534]=64;
sine[1535]=64;
sine[1536]=64;
sine[1537]=64;
sine[1538]=64;
sine[1539]=64;
sine[1540]=64;
sine[1541]=64;
sine[1542]=64;
sine[1543]=64;
sine[1544]=64;
sine[1545]=64;
sine[1546]=65;
sine[1547]=65;
sine[1548]=65;
sine[1549]=65;
sine[1550]=65;
sine[1551]=65;
sine[1552]=65;
sine[1553]=65;
sine[1554]=65;
sine[1555]=65;
sine[1556]=65;
sine[1557]=65;
sine[1558]=65;
sine[1559]=65;
sine[1560]=65;
sine[1561]=65;
sine[1562]=65;
sine[1563]=65;
sine[1564]=65;
sine[1565]=65;
sine[1566]=65;
sine[1567]=65;
sine[1568]=65;
sine[1569]=65;
sine[1570]=65;
sine[1571]=65;
sine[1572]=65;
sine[1573]=65;
sine[1574]=65;
sine[1575]=65;
sine[1576]=65;
sine[1577]=65;
sine[1578]=65;
sine[1579]=65;
sine[1580]=65;
sine[1581]=65;
sine[1582]=65;
sine[1583]=66;
sine[1584]=66;
sine[1585]=66;
sine[1586]=66;
sine[1587]=66;
sine[1588]=66;
sine[1589]=66;
sine[1590]=66;
sine[1591]=66;
sine[1592]=66;
sine[1593]=66;
sine[1594]=66;
sine[1595]=66;
sine[1596]=66;
sine[1597]=66;
sine[1598]=66;
sine[1599]=66;
sine[1600]=66;
sine[1601]=66;
sine[1602]=66;
sine[1603]=66;
sine[1604]=66;
sine[1605]=66;
sine[1606]=66;
sine[1607]=66;
sine[1608]=66;
sine[1609]=66;
sine[1610]=66;
sine[1611]=66;
sine[1612]=66;
sine[1613]=66;
sine[1614]=66;
sine[1615]=66;
sine[1616]=66;
sine[1617]=66;
sine[1618]=66;
sine[1619]=66;
sine[1620]=66;
sine[1621]=67;
sine[1622]=67;
sine[1623]=67;
sine[1624]=67;
sine[1625]=67;
sine[1626]=67;
sine[1627]=67;
sine[1628]=67;
sine[1629]=67;
sine[1630]=67;
sine[1631]=67;
sine[1632]=67;
sine[1633]=67;
sine[1634]=67;
sine[1635]=67;
sine[1636]=67;
sine[1637]=67;
sine[1638]=67;
sine[1639]=67;
sine[1640]=67;
sine[1641]=67;
sine[1642]=67;
sine[1643]=67;
sine[1644]=67;
sine[1645]=67;
sine[1646]=67;
sine[1647]=67;
sine[1648]=67;
sine[1649]=67;
sine[1650]=67;
sine[1651]=67;
sine[1652]=67;
sine[1653]=67;
sine[1654]=67;
sine[1655]=67;
sine[1656]=67;
sine[1657]=67;
sine[1658]=67;
sine[1659]=67;
sine[1660]=67;
sine[1661]=68;
sine[1662]=68;
sine[1663]=68;
sine[1664]=68;
sine[1665]=68;
sine[1666]=68;
sine[1667]=68;
sine[1668]=68;
sine[1669]=68;
sine[1670]=68;
sine[1671]=68;
sine[1672]=68;
sine[1673]=68;
sine[1674]=68;
sine[1675]=68;
sine[1676]=68;
sine[1677]=68;
sine[1678]=68;
sine[1679]=68;
sine[1680]=68;
sine[1681]=68;
sine[1682]=68;
sine[1683]=68;
sine[1684]=68;
sine[1685]=68;
sine[1686]=68;
sine[1687]=68;
sine[1688]=68;
sine[1689]=68;
sine[1690]=68;
sine[1691]=68;
sine[1692]=68;
sine[1693]=68;
sine[1694]=68;
sine[1695]=68;
sine[1696]=68;
sine[1697]=68;
sine[1698]=68;
sine[1699]=68;
sine[1700]=68;
sine[1701]=68;
sine[1702]=69;
sine[1703]=69;
sine[1704]=69;
sine[1705]=69;
sine[1706]=69;
sine[1707]=69;
sine[1708]=69;
sine[1709]=69;
sine[1710]=69;
sine[1711]=69;
sine[1712]=69;
sine[1713]=69;
sine[1714]=69;
sine[1715]=69;
sine[1716]=69;
sine[1717]=69;
sine[1718]=69;
sine[1719]=69;
sine[1720]=69;
sine[1721]=69;
sine[1722]=69;
sine[1723]=69;
sine[1724]=69;
sine[1725]=69;
sine[1726]=69;
sine[1727]=69;
sine[1728]=69;
sine[1729]=69;
sine[1730]=69;
sine[1731]=69;
sine[1732]=69;
sine[1733]=69;
sine[1734]=69;
sine[1735]=69;
sine[1736]=69;
sine[1737]=69;
sine[1738]=69;
sine[1739]=69;
sine[1740]=69;
sine[1741]=69;
sine[1742]=69;
sine[1743]=69;
sine[1744]=69;
sine[1745]=69;
sine[1746]=70;
sine[1747]=70;
sine[1748]=70;
sine[1749]=70;
sine[1750]=70;
sine[1751]=70;
sine[1752]=70;
sine[1753]=70;
sine[1754]=70;
sine[1755]=70;
sine[1756]=70;
sine[1757]=70;
sine[1758]=70;
sine[1759]=70;
sine[1760]=70;
sine[1761]=70;
sine[1762]=70;
sine[1763]=70;
sine[1764]=70;
sine[1765]=70;
sine[1766]=70;
sine[1767]=70;
sine[1768]=70;
sine[1769]=70;
sine[1770]=70;
sine[1771]=70;
sine[1772]=70;
sine[1773]=70;
sine[1774]=70;
sine[1775]=70;
sine[1776]=70;
sine[1777]=70;
sine[1778]=70;
sine[1779]=70;
sine[1780]=70;
sine[1781]=70;
sine[1782]=70;
sine[1783]=70;
sine[1784]=70;
sine[1785]=70;
sine[1786]=70;
sine[1787]=70;
sine[1788]=70;
sine[1789]=70;
sine[1790]=70;
sine[1791]=71;
sine[1792]=71;
sine[1793]=71;
sine[1794]=71;
sine[1795]=71;
sine[1796]=71;
sine[1797]=71;
sine[1798]=71;
sine[1799]=71;
sine[1800]=71;
sine[1801]=71;
sine[1802]=71;
sine[1803]=71;
sine[1804]=71;
sine[1805]=71;
sine[1806]=71;
sine[1807]=71;
sine[1808]=71;
sine[1809]=71;
sine[1810]=71;
sine[1811]=71;
sine[1812]=71;
sine[1813]=71;
sine[1814]=71;
sine[1815]=71;
sine[1816]=71;
sine[1817]=71;
sine[1818]=71;
sine[1819]=71;
sine[1820]=71;
sine[1821]=71;
sine[1822]=71;
sine[1823]=71;
sine[1824]=71;
sine[1825]=71;
sine[1826]=71;
sine[1827]=71;
sine[1828]=71;
sine[1829]=71;
sine[1830]=71;
sine[1831]=71;
sine[1832]=71;
sine[1833]=71;
sine[1834]=71;
sine[1835]=71;
sine[1836]=71;
sine[1837]=71;
sine[1838]=71;
sine[1839]=71;
sine[1840]=72;
sine[1841]=72;
sine[1842]=72;
sine[1843]=72;
sine[1844]=72;
sine[1845]=72;
sine[1846]=72;
sine[1847]=72;
sine[1848]=72;
sine[1849]=72;
sine[1850]=72;
sine[1851]=72;
sine[1852]=72;
sine[1853]=72;
sine[1854]=72;
sine[1855]=72;
sine[1856]=72;
sine[1857]=72;
sine[1858]=72;
sine[1859]=72;
sine[1860]=72;
sine[1861]=72;
sine[1862]=72;
sine[1863]=72;
sine[1864]=72;
sine[1865]=72;
sine[1866]=72;
sine[1867]=72;
sine[1868]=72;
sine[1869]=72;
sine[1870]=72;
sine[1871]=72;
sine[1872]=72;
sine[1873]=72;
sine[1874]=72;
sine[1875]=72;
sine[1876]=72;
sine[1877]=72;
sine[1878]=72;
sine[1879]=72;
sine[1880]=72;
sine[1881]=72;
sine[1882]=72;
sine[1883]=72;
sine[1884]=72;
sine[1885]=72;
sine[1886]=72;
sine[1887]=72;
sine[1888]=72;
sine[1889]=72;
sine[1890]=72;
sine[1891]=72;
sine[1892]=72;
sine[1893]=73;
sine[1894]=73;
sine[1895]=73;
sine[1896]=73;
sine[1897]=73;
sine[1898]=73;
sine[1899]=73;
sine[1900]=73;
sine[1901]=73;
sine[1902]=73;
sine[1903]=73;
sine[1904]=73;
sine[1905]=73;
sine[1906]=73;
sine[1907]=73;
sine[1908]=73;
sine[1909]=73;
sine[1910]=73;
sine[1911]=73;
sine[1912]=73;
sine[1913]=73;
sine[1914]=73;
sine[1915]=73;
sine[1916]=73;
sine[1917]=73;
sine[1918]=73;
sine[1919]=73;
sine[1920]=73;
sine[1921]=73;
sine[1922]=73;
sine[1923]=73;
sine[1924]=73;
sine[1925]=73;
sine[1926]=73;
sine[1927]=73;
sine[1928]=73;
sine[1929]=73;
sine[1930]=73;
sine[1931]=73;
sine[1932]=73;
sine[1933]=73;
sine[1934]=73;
sine[1935]=73;
sine[1936]=73;
sine[1937]=73;
sine[1938]=73;
sine[1939]=73;
sine[1940]=73;
sine[1941]=73;
sine[1942]=73;
sine[1943]=73;
sine[1944]=73;
sine[1945]=73;
sine[1946]=73;
sine[1947]=73;
sine[1948]=73;
sine[1949]=73;
sine[1950]=74;
sine[1951]=74;
sine[1952]=74;
sine[1953]=74;
sine[1954]=74;
sine[1955]=74;
sine[1956]=74;
sine[1957]=74;
sine[1958]=74;
sine[1959]=74;
sine[1960]=74;
sine[1961]=74;
sine[1962]=74;
sine[1963]=74;
sine[1964]=74;
sine[1965]=74;
sine[1966]=74;
sine[1967]=74;
sine[1968]=74;
sine[1969]=74;
sine[1970]=74;
sine[1971]=74;
sine[1972]=74;
sine[1973]=74;
sine[1974]=74;
sine[1975]=74;
sine[1976]=74;
sine[1977]=74;
sine[1978]=74;
sine[1979]=74;
sine[1980]=74;
sine[1981]=74;
sine[1982]=74;
sine[1983]=74;
sine[1984]=74;
sine[1985]=74;
sine[1986]=74;
sine[1987]=74;
sine[1988]=74;
sine[1989]=74;
sine[1990]=74;
sine[1991]=74;
sine[1992]=74;
sine[1993]=74;
sine[1994]=74;
sine[1995]=74;
sine[1996]=74;
sine[1997]=74;
sine[1998]=74;
sine[1999]=74;
sine[2000]=74;
sine[2001]=74;
sine[2002]=74;
sine[2003]=74;
sine[2004]=74;
sine[2005]=74;
sine[2006]=74;
sine[2007]=74;
sine[2008]=74;
sine[2009]=74;
sine[2010]=74;
sine[2011]=74;
sine[2012]=74;
sine[2013]=74;
sine[2014]=75;
sine[2015]=75;
sine[2016]=75;
sine[2017]=75;
sine[2018]=75;
sine[2019]=75;
sine[2020]=75;
sine[2021]=75;
sine[2022]=75;
sine[2023]=75;
sine[2024]=75;
sine[2025]=75;
sine[2026]=75;
sine[2027]=75;
sine[2028]=75;
sine[2029]=75;
sine[2030]=75;
sine[2031]=75;
sine[2032]=75;
sine[2033]=75;
sine[2034]=75;
sine[2035]=75;
sine[2036]=75;
sine[2037]=75;
sine[2038]=75;
sine[2039]=75;
sine[2040]=75;
sine[2041]=75;
sine[2042]=75;
sine[2043]=75;
sine[2044]=75;
sine[2045]=75;
sine[2046]=75;
sine[2047]=75;
sine[2048]=75;
sine[2049]=75;
sine[2050]=75;
sine[2051]=75;
sine[2052]=75;
sine[2053]=75;
sine[2054]=75;
sine[2055]=75;
sine[2056]=75;
sine[2057]=75;
sine[2058]=75;
sine[2059]=75;
sine[2060]=75;
sine[2061]=75;
sine[2062]=75;
sine[2063]=75;
sine[2064]=75;
sine[2065]=75;
sine[2066]=75;
sine[2067]=75;
sine[2068]=75;
sine[2069]=75;
sine[2070]=75;
sine[2071]=75;
sine[2072]=75;
sine[2073]=75;
sine[2074]=75;
sine[2075]=75;
sine[2076]=75;
sine[2077]=75;
sine[2078]=75;
sine[2079]=75;
sine[2080]=75;
sine[2081]=75;
sine[2082]=75;
sine[2083]=75;
sine[2084]=75;
sine[2085]=75;
sine[2086]=75;
sine[2087]=76;
sine[2088]=76;
sine[2089]=76;
sine[2090]=76;
sine[2091]=76;
sine[2092]=76;
sine[2093]=76;
sine[2094]=76;
sine[2095]=76;
sine[2096]=76;
sine[2097]=76;
sine[2098]=76;
sine[2099]=76;
sine[2100]=76;
sine[2101]=76;
sine[2102]=76;
sine[2103]=76;
sine[2104]=76;
sine[2105]=76;
sine[2106]=76;
sine[2107]=76;
sine[2108]=76;
sine[2109]=76;
sine[2110]=76;
sine[2111]=76;
sine[2112]=76;
sine[2113]=76;
sine[2114]=76;
sine[2115]=76;
sine[2116]=76;
sine[2117]=76;
sine[2118]=76;
sine[2119]=76;
sine[2120]=76;
sine[2121]=76;
sine[2122]=76;
sine[2123]=76;
sine[2124]=76;
sine[2125]=76;
sine[2126]=76;
sine[2127]=76;
sine[2128]=76;
sine[2129]=76;
sine[2130]=76;
sine[2131]=76;
sine[2132]=76;
sine[2133]=76;
sine[2134]=76;
sine[2135]=76;
sine[2136]=76;
sine[2137]=76;
sine[2138]=76;
sine[2139]=76;
sine[2140]=76;
sine[2141]=76;
sine[2142]=76;
sine[2143]=76;
sine[2144]=76;
sine[2145]=76;
sine[2146]=76;
sine[2147]=76;
sine[2148]=76;
sine[2149]=76;
sine[2150]=76;
sine[2151]=76;
sine[2152]=76;
sine[2153]=76;
sine[2154]=76;
sine[2155]=76;
sine[2156]=76;
sine[2157]=76;
sine[2158]=76;
sine[2159]=76;
sine[2160]=76;
sine[2161]=76;
sine[2162]=76;
sine[2163]=76;
sine[2164]=76;
sine[2165]=76;
sine[2166]=76;
sine[2167]=76;
sine[2168]=76;
sine[2169]=76;
sine[2170]=76;
sine[2171]=76;
sine[2172]=76;
sine[2173]=76;
sine[2174]=76;
sine[2175]=77;
sine[2176]=77;
sine[2177]=77;
sine[2178]=77;
sine[2179]=77;
sine[2180]=77;
sine[2181]=77;
sine[2182]=77;
sine[2183]=77;
sine[2184]=77;
sine[2185]=77;
sine[2186]=77;
sine[2187]=77;
sine[2188]=77;
sine[2189]=77;
sine[2190]=77;
sine[2191]=77;
sine[2192]=77;
sine[2193]=77;
sine[2194]=77;
sine[2195]=77;
sine[2196]=77;
sine[2197]=77;
sine[2198]=77;
sine[2199]=77;
sine[2200]=77;
sine[2201]=77;
sine[2202]=77;
sine[2203]=77;
sine[2204]=77;
sine[2205]=77;
sine[2206]=77;
sine[2207]=77;
sine[2208]=77;
sine[2209]=77;
sine[2210]=77;
sine[2211]=77;
sine[2212]=77;
sine[2213]=77;
sine[2214]=77;
sine[2215]=77;
sine[2216]=77;
sine[2217]=77;
sine[2218]=77;
sine[2219]=77;
sine[2220]=77;
sine[2221]=77;
sine[2222]=77;
sine[2223]=77;
sine[2224]=77;
sine[2225]=77;
sine[2226]=77;
sine[2227]=77;
sine[2228]=77;
sine[2229]=77;
sine[2230]=77;
sine[2231]=77;
sine[2232]=77;
sine[2233]=77;
sine[2234]=77;
sine[2235]=77;
sine[2236]=77;
sine[2237]=77;
sine[2238]=77;
sine[2239]=77;
sine[2240]=77;
sine[2241]=77;
sine[2242]=77;
sine[2243]=77;
sine[2244]=77;
sine[2245]=77;
sine[2246]=77;
sine[2247]=77;
sine[2248]=77;
sine[2249]=77;
sine[2250]=77;
sine[2251]=77;
sine[2252]=77;
sine[2253]=77;
sine[2254]=77;
sine[2255]=77;
sine[2256]=77;
sine[2257]=77;
sine[2258]=77;
sine[2259]=77;
sine[2260]=77;
sine[2261]=77;
sine[2262]=77;
sine[2263]=77;
sine[2264]=77;
sine[2265]=77;
sine[2266]=77;
sine[2267]=77;
sine[2268]=77;
sine[2269]=77;
sine[2270]=77;
sine[2271]=77;
sine[2272]=77;
sine[2273]=77;
sine[2274]=77;
sine[2275]=77;
sine[2276]=77;
sine[2277]=77;
sine[2278]=77;
sine[2279]=77;
sine[2280]=77;
sine[2281]=77;
sine[2282]=77;
sine[2283]=77;
sine[2284]=77;
sine[2285]=77;
sine[2286]=77;
sine[2287]=77;
sine[2288]=77;
sine[2289]=77;
sine[2290]=77;
sine[2291]=77;
sine[2292]=77;
sine[2293]=77;
sine[2294]=77;
sine[2295]=77;
sine[2296]=77;
sine[2297]=77;
sine[2298]=77;
sine[2299]=78;
sine[2300]=78;
sine[2301]=78;
sine[2302]=78;
sine[2303]=78;
sine[2304]=78;
sine[2305]=78;
sine[2306]=78;
sine[2307]=78;
sine[2308]=78;
sine[2309]=78;
sine[2310]=78;
sine[2311]=78;
sine[2312]=78;
sine[2313]=78;
sine[2314]=78;
sine[2315]=78;
sine[2316]=78;
sine[2317]=78;
sine[2318]=78;
sine[2319]=78;
sine[2320]=78;
sine[2321]=78;
sine[2322]=78;
sine[2323]=78;
sine[2324]=78;
sine[2325]=78;
sine[2326]=78;
sine[2327]=78;
sine[2328]=78;
sine[2329]=78;
sine[2330]=78;
sine[2331]=78;
sine[2332]=78;
sine[2333]=78;
sine[2334]=78;
sine[2335]=78;
sine[2336]=78;
sine[2337]=78;
sine[2338]=78;
sine[2339]=78;
sine[2340]=78;
sine[2341]=78;
sine[2342]=78;
sine[2343]=78;
sine[2344]=78;
sine[2345]=78;
sine[2346]=78;
sine[2347]=78;
sine[2348]=78;
sine[2349]=78;
sine[2350]=78;
sine[2351]=78;
sine[2352]=78;
sine[2353]=78;
sine[2354]=78;
sine[2355]=78;
sine[2356]=78;
sine[2357]=78;
sine[2358]=78;
sine[2359]=78;
sine[2360]=78;
sine[2361]=78;
sine[2362]=78;
sine[2363]=78;
sine[2364]=78;
sine[2365]=78;
sine[2366]=78;
sine[2367]=78;
sine[2368]=78;
sine[2369]=78;
sine[2370]=78;
sine[2371]=78;
sine[2372]=78;
sine[2373]=78;
sine[2374]=78;
sine[2375]=78;
sine[2376]=78;
sine[2377]=78;
sine[2378]=78;
sine[2379]=78;
sine[2380]=78;
sine[2381]=78;
sine[2382]=78;
sine[2383]=78;
sine[2384]=78;
sine[2385]=78;
sine[2386]=78;
sine[2387]=78;
sine[2388]=78;
sine[2389]=78;
sine[2390]=78;
sine[2391]=78;
sine[2392]=78;
sine[2393]=78;
sine[2394]=78;
sine[2395]=78;
sine[2396]=78;
sine[2397]=78;
sine[2398]=78;
sine[2399]=78;
sine[2400]=78;
sine[2401]=78;
sine[2402]=78;
sine[2403]=78;
sine[2404]=78;
sine[2405]=78;
sine[2406]=78;
sine[2407]=78;
sine[2408]=78;
sine[2409]=78;
sine[2410]=78;
sine[2411]=78;
sine[2412]=78;
sine[2413]=78;
sine[2414]=78;
sine[2415]=78;
sine[2416]=78;
sine[2417]=78;
sine[2418]=78;
sine[2419]=78;
sine[2420]=78;
sine[2421]=78;
sine[2422]=78;
sine[2423]=78;
sine[2424]=78;
sine[2425]=78;
sine[2426]=78;
sine[2427]=78;
sine[2428]=78;
sine[2429]=78;
sine[2430]=78;
sine[2431]=78;
sine[2432]=78;
sine[2433]=78;
sine[2434]=78;
sine[2435]=78;
sine[2436]=78;
sine[2437]=78;
sine[2438]=78;
sine[2439]=78;
sine[2440]=78;
sine[2441]=78;
sine[2442]=78;
sine[2443]=78;
sine[2444]=78;
sine[2445]=78;
sine[2446]=78;
sine[2447]=78;
sine[2448]=78;
sine[2449]=78;
sine[2450]=78;
sine[2451]=78;
sine[2452]=78;
sine[2453]=78;
sine[2454]=78;
sine[2455]=78;
sine[2456]=78;
sine[2457]=78;
sine[2458]=78;
sine[2459]=78;
sine[2460]=78;
sine[2461]=78;
sine[2462]=78;
sine[2463]=78;
sine[2464]=78;
sine[2465]=78;
sine[2466]=78;
sine[2467]=78;
sine[2468]=78;
sine[2469]=78;
sine[2470]=78;
sine[2471]=78;
sine[2472]=78;
sine[2473]=78;
sine[2474]=78;
sine[2475]=78;
sine[2476]=78;
sine[2477]=78;
sine[2478]=78;
sine[2479]=78;
sine[2480]=78;
sine[2481]=78;
sine[2482]=78;
sine[2483]=78;
sine[2484]=78;
sine[2485]=78;
sine[2486]=78;
sine[2487]=78;
sine[2488]=78;
sine[2489]=78;
sine[2490]=78;
sine[2491]=78;
sine[2492]=78;
sine[2493]=78;
sine[2494]=78;
sine[2495]=78;
sine[2496]=78;
sine[2497]=78;
sine[2498]=78;
sine[2499]=78;
sine[2500]=78;
sine[2501]=78;
sine[2502]=78;
sine[2503]=78;
sine[2504]=78;
sine[2505]=78;
sine[2506]=78;
sine[2507]=78;
sine[2508]=78;
sine[2509]=78;
sine[2510]=78;
sine[2511]=78;
sine[2512]=78;
sine[2513]=78;
sine[2514]=78;
sine[2515]=78;
sine[2516]=78;
sine[2517]=78;
sine[2518]=78;
sine[2519]=78;
sine[2520]=78;
sine[2521]=78;
sine[2522]=78;
sine[2523]=78;
sine[2524]=78;
sine[2525]=78;
sine[2526]=78;
sine[2527]=78;
sine[2528]=78;
sine[2529]=78;
sine[2530]=78;
sine[2531]=78;
sine[2532]=78;
sine[2533]=78;
sine[2534]=78;
sine[2535]=78;
sine[2536]=78;
sine[2537]=78;
sine[2538]=78;
sine[2539]=78;
sine[2540]=78;
sine[2541]=78;
sine[2542]=78;
sine[2543]=78;
sine[2544]=78;
sine[2545]=78;
sine[2546]=78;
sine[2547]=78;
sine[2548]=78;
sine[2549]=78;
sine[2550]=78;
sine[2551]=78;
sine[2552]=78;
sine[2553]=78;
sine[2554]=78;
sine[2555]=78;
sine[2556]=78;
sine[2557]=78;
sine[2558]=78;
sine[2559]=78;
sine[2560]=78;
sine[2561]=78;
sine[2562]=78;
sine[2563]=78;
sine[2564]=78;
sine[2565]=78;
sine[2566]=78;
sine[2567]=78;
sine[2568]=78;
sine[2569]=78;
sine[2570]=78;
sine[2571]=78;
sine[2572]=78;
sine[2573]=78;
sine[2574]=78;
sine[2575]=78;
sine[2576]=78;
sine[2577]=78;
sine[2578]=78;
sine[2579]=78;
sine[2580]=78;
sine[2581]=78;
sine[2582]=78;
sine[2583]=78;
sine[2584]=78;
sine[2585]=78;
sine[2586]=78;
sine[2587]=78;
sine[2588]=78;
sine[2589]=78;
sine[2590]=78;
sine[2591]=78;
sine[2592]=78;
sine[2593]=78;
sine[2594]=78;
sine[2595]=78;
sine[2596]=78;
sine[2597]=78;
sine[2598]=78;
sine[2599]=78;
sine[2600]=78;
sine[2601]=78;
sine[2602]=78;
sine[2603]=78;
sine[2604]=78;
sine[2605]=78;
sine[2606]=78;
sine[2607]=78;
sine[2608]=78;
sine[2609]=78;
sine[2610]=78;
sine[2611]=78;
sine[2612]=78;
sine[2613]=78;
sine[2614]=78;
sine[2615]=78;
sine[2616]=78;
sine[2617]=78;
sine[2618]=78;
sine[2619]=78;
sine[2620]=78;
sine[2621]=78;
sine[2622]=78;
sine[2623]=78;
sine[2624]=78;
sine[2625]=78;
sine[2626]=78;
sine[2627]=78;
sine[2628]=78;
sine[2629]=78;
sine[2630]=78;
sine[2631]=78;
sine[2632]=78;
sine[2633]=78;
sine[2634]=78;
sine[2635]=78;
sine[2636]=78;
sine[2637]=78;
sine[2638]=78;
sine[2639]=78;
sine[2640]=78;
sine[2641]=78;
sine[2642]=78;
sine[2643]=78;
sine[2644]=78;
sine[2645]=78;
sine[2646]=78;
sine[2647]=78;
sine[2648]=78;
sine[2649]=78;
sine[2650]=78;
sine[2651]=78;
sine[2652]=78;
sine[2653]=78;
sine[2654]=78;
sine[2655]=78;
sine[2656]=78;
sine[2657]=78;
sine[2658]=78;
sine[2659]=78;
sine[2660]=78;
sine[2661]=78;
sine[2662]=78;
sine[2663]=78;
sine[2664]=78;
sine[2665]=78;
sine[2666]=78;
sine[2667]=78;
sine[2668]=78;
sine[2669]=78;
sine[2670]=78;
sine[2671]=78;
sine[2672]=78;
sine[2673]=78;
sine[2674]=78;
sine[2675]=78;
sine[2676]=78;
sine[2677]=78;
sine[2678]=78;
sine[2679]=78;
sine[2680]=78;
sine[2681]=78;
sine[2682]=78;
sine[2683]=78;
sine[2684]=78;
sine[2685]=78;
sine[2686]=78;
sine[2687]=78;
sine[2688]=78;
sine[2689]=78;
sine[2690]=78;
sine[2691]=78;
sine[2692]=78;
sine[2693]=78;
sine[2694]=78;
sine[2695]=78;
sine[2696]=78;
sine[2697]=78;
sine[2698]=78;
sine[2699]=78;
sine[2700]=78;
sine[2701]=78;
sine[2702]=77;
sine[2703]=77;
sine[2704]=77;
sine[2705]=77;
sine[2706]=77;
sine[2707]=77;
sine[2708]=77;
sine[2709]=77;
sine[2710]=77;
sine[2711]=77;
sine[2712]=77;
sine[2713]=77;
sine[2714]=77;
sine[2715]=77;
sine[2716]=77;
sine[2717]=77;
sine[2718]=77;
sine[2719]=77;
sine[2720]=77;
sine[2721]=77;
sine[2722]=77;
sine[2723]=77;
sine[2724]=77;
sine[2725]=77;
sine[2726]=77;
sine[2727]=77;
sine[2728]=77;
sine[2729]=77;
sine[2730]=77;
sine[2731]=77;
sine[2732]=77;
sine[2733]=77;
sine[2734]=77;
sine[2735]=77;
sine[2736]=77;
sine[2737]=77;
sine[2738]=77;
sine[2739]=77;
sine[2740]=77;
sine[2741]=77;
sine[2742]=77;
sine[2743]=77;
sine[2744]=77;
sine[2745]=77;
sine[2746]=77;
sine[2747]=77;
sine[2748]=77;
sine[2749]=77;
sine[2750]=77;
sine[2751]=77;
sine[2752]=77;
sine[2753]=77;
sine[2754]=77;
sine[2755]=77;
sine[2756]=77;
sine[2757]=77;
sine[2758]=77;
sine[2759]=77;
sine[2760]=77;
sine[2761]=77;
sine[2762]=77;
sine[2763]=77;
sine[2764]=77;
sine[2765]=77;
sine[2766]=77;
sine[2767]=77;
sine[2768]=77;
sine[2769]=77;
sine[2770]=77;
sine[2771]=77;
sine[2772]=77;
sine[2773]=77;
sine[2774]=77;
sine[2775]=77;
sine[2776]=77;
sine[2777]=77;
sine[2778]=77;
sine[2779]=77;
sine[2780]=77;
sine[2781]=77;
sine[2782]=77;
sine[2783]=77;
sine[2784]=77;
sine[2785]=77;
sine[2786]=77;
sine[2787]=77;
sine[2788]=77;
sine[2789]=77;
sine[2790]=77;
sine[2791]=77;
sine[2792]=77;
sine[2793]=77;
sine[2794]=77;
sine[2795]=77;
sine[2796]=77;
sine[2797]=77;
sine[2798]=77;
sine[2799]=77;
sine[2800]=77;
sine[2801]=77;
sine[2802]=77;
sine[2803]=77;
sine[2804]=77;
sine[2805]=77;
sine[2806]=77;
sine[2807]=77;
sine[2808]=77;
sine[2809]=77;
sine[2810]=77;
sine[2811]=77;
sine[2812]=77;
sine[2813]=77;
sine[2814]=77;
sine[2815]=77;
sine[2816]=77;
sine[2817]=77;
sine[2818]=77;
sine[2819]=77;
sine[2820]=77;
sine[2821]=77;
sine[2822]=77;
sine[2823]=77;
sine[2824]=77;
sine[2825]=77;
sine[2826]=76;
sine[2827]=76;
sine[2828]=76;
sine[2829]=76;
sine[2830]=76;
sine[2831]=76;
sine[2832]=76;
sine[2833]=76;
sine[2834]=76;
sine[2835]=76;
sine[2836]=76;
sine[2837]=76;
sine[2838]=76;
sine[2839]=76;
sine[2840]=76;
sine[2841]=76;
sine[2842]=76;
sine[2843]=76;
sine[2844]=76;
sine[2845]=76;
sine[2846]=76;
sine[2847]=76;
sine[2848]=76;
sine[2849]=76;
sine[2850]=76;
sine[2851]=76;
sine[2852]=76;
sine[2853]=76;
sine[2854]=76;
sine[2855]=76;
sine[2856]=76;
sine[2857]=76;
sine[2858]=76;
sine[2859]=76;
sine[2860]=76;
sine[2861]=76;
sine[2862]=76;
sine[2863]=76;
sine[2864]=76;
sine[2865]=76;
sine[2866]=76;
sine[2867]=76;
sine[2868]=76;
sine[2869]=76;
sine[2870]=76;
sine[2871]=76;
sine[2872]=76;
sine[2873]=76;
sine[2874]=76;
sine[2875]=76;
sine[2876]=76;
sine[2877]=76;
sine[2878]=76;
sine[2879]=76;
sine[2880]=76;
sine[2881]=76;
sine[2882]=76;
sine[2883]=76;
sine[2884]=76;
sine[2885]=76;
sine[2886]=76;
sine[2887]=76;
sine[2888]=76;
sine[2889]=76;
sine[2890]=76;
sine[2891]=76;
sine[2892]=76;
sine[2893]=76;
sine[2894]=76;
sine[2895]=76;
sine[2896]=76;
sine[2897]=76;
sine[2898]=76;
sine[2899]=76;
sine[2900]=76;
sine[2901]=76;
sine[2902]=76;
sine[2903]=76;
sine[2904]=76;
sine[2905]=76;
sine[2906]=76;
sine[2907]=76;
sine[2908]=76;
sine[2909]=76;
sine[2910]=76;
sine[2911]=76;
sine[2912]=76;
sine[2913]=76;
sine[2914]=75;
sine[2915]=75;
sine[2916]=75;
sine[2917]=75;
sine[2918]=75;
sine[2919]=75;
sine[2920]=75;
sine[2921]=75;
sine[2922]=75;
sine[2923]=75;
sine[2924]=75;
sine[2925]=75;
sine[2926]=75;
sine[2927]=75;
sine[2928]=75;
sine[2929]=75;
sine[2930]=75;
sine[2931]=75;
sine[2932]=75;
sine[2933]=75;
sine[2934]=75;
sine[2935]=75;
sine[2936]=75;
sine[2937]=75;
sine[2938]=75;
sine[2939]=75;
sine[2940]=75;
sine[2941]=75;
sine[2942]=75;
sine[2943]=75;
sine[2944]=75;
sine[2945]=75;
sine[2946]=75;
sine[2947]=75;
sine[2948]=75;
sine[2949]=75;
sine[2950]=75;
sine[2951]=75;
sine[2952]=75;
sine[2953]=75;
sine[2954]=75;
sine[2955]=75;
sine[2956]=75;
sine[2957]=75;
sine[2958]=75;
sine[2959]=75;
sine[2960]=75;
sine[2961]=75;
sine[2962]=75;
sine[2963]=75;
sine[2964]=75;
sine[2965]=75;
sine[2966]=75;
sine[2967]=75;
sine[2968]=75;
sine[2969]=75;
sine[2970]=75;
sine[2971]=75;
sine[2972]=75;
sine[2973]=75;
sine[2974]=75;
sine[2975]=75;
sine[2976]=75;
sine[2977]=75;
sine[2978]=75;
sine[2979]=75;
sine[2980]=75;
sine[2981]=75;
sine[2982]=75;
sine[2983]=75;
sine[2984]=75;
sine[2985]=75;
sine[2986]=75;
sine[2987]=74;
sine[2988]=74;
sine[2989]=74;
sine[2990]=74;
sine[2991]=74;
sine[2992]=74;
sine[2993]=74;
sine[2994]=74;
sine[2995]=74;
sine[2996]=74;
sine[2997]=74;
sine[2998]=74;
sine[2999]=74;
sine[3000]=74;
sine[3001]=74;
sine[3002]=74;
sine[3003]=74;
sine[3004]=74;
sine[3005]=74;
sine[3006]=74;
sine[3007]=74;
sine[3008]=74;
sine[3009]=74;
sine[3010]=74;
sine[3011]=74;
sine[3012]=74;
sine[3013]=74;
sine[3014]=74;
sine[3015]=74;
sine[3016]=74;
sine[3017]=74;
sine[3018]=74;
sine[3019]=74;
sine[3020]=74;
sine[3021]=74;
sine[3022]=74;
sine[3023]=74;
sine[3024]=74;
sine[3025]=74;
sine[3026]=74;
sine[3027]=74;
sine[3028]=74;
sine[3029]=74;
sine[3030]=74;
sine[3031]=74;
sine[3032]=74;
sine[3033]=74;
sine[3034]=74;
sine[3035]=74;
sine[3036]=74;
sine[3037]=74;
sine[3038]=74;
sine[3039]=74;
sine[3040]=74;
sine[3041]=74;
sine[3042]=74;
sine[3043]=74;
sine[3044]=74;
sine[3045]=74;
sine[3046]=74;
sine[3047]=74;
sine[3048]=74;
sine[3049]=74;
sine[3050]=74;
sine[3051]=73;
sine[3052]=73;
sine[3053]=73;
sine[3054]=73;
sine[3055]=73;
sine[3056]=73;
sine[3057]=73;
sine[3058]=73;
sine[3059]=73;
sine[3060]=73;
sine[3061]=73;
sine[3062]=73;
sine[3063]=73;
sine[3064]=73;
sine[3065]=73;
sine[3066]=73;
sine[3067]=73;
sine[3068]=73;
sine[3069]=73;
sine[3070]=73;
sine[3071]=73;
sine[3072]=73;
sine[3073]=73;
sine[3074]=73;
sine[3075]=73;
sine[3076]=73;
sine[3077]=73;
sine[3078]=73;
sine[3079]=73;
sine[3080]=73;
sine[3081]=73;
sine[3082]=73;
sine[3083]=73;
sine[3084]=73;
sine[3085]=73;
sine[3086]=73;
sine[3087]=73;
sine[3088]=73;
sine[3089]=73;
sine[3090]=73;
sine[3091]=73;
sine[3092]=73;
sine[3093]=73;
sine[3094]=73;
sine[3095]=73;
sine[3096]=73;
sine[3097]=73;
sine[3098]=73;
sine[3099]=73;
sine[3100]=73;
sine[3101]=73;
sine[3102]=73;
sine[3103]=73;
sine[3104]=73;
sine[3105]=73;
sine[3106]=73;
sine[3107]=73;
sine[3108]=72;
sine[3109]=72;
sine[3110]=72;
sine[3111]=72;
sine[3112]=72;
sine[3113]=72;
sine[3114]=72;
sine[3115]=72;
sine[3116]=72;
sine[3117]=72;
sine[3118]=72;
sine[3119]=72;
sine[3120]=72;
sine[3121]=72;
sine[3122]=72;
sine[3123]=72;
sine[3124]=72;
sine[3125]=72;
sine[3126]=72;
sine[3127]=72;
sine[3128]=72;
sine[3129]=72;
sine[3130]=72;
sine[3131]=72;
sine[3132]=72;
sine[3133]=72;
sine[3134]=72;
sine[3135]=72;
sine[3136]=72;
sine[3137]=72;
sine[3138]=72;
sine[3139]=72;
sine[3140]=72;
sine[3141]=72;
sine[3142]=72;
sine[3143]=72;
sine[3144]=72;
sine[3145]=72;
sine[3146]=72;
sine[3147]=72;
sine[3148]=72;
sine[3149]=72;
sine[3150]=72;
sine[3151]=72;
sine[3152]=72;
sine[3153]=72;
sine[3154]=72;
sine[3155]=72;
sine[3156]=72;
sine[3157]=72;
sine[3158]=72;
sine[3159]=72;
sine[3160]=72;
sine[3161]=71;
sine[3162]=71;
sine[3163]=71;
sine[3164]=71;
sine[3165]=71;
sine[3166]=71;
sine[3167]=71;
sine[3168]=71;
sine[3169]=71;
sine[3170]=71;
sine[3171]=71;
sine[3172]=71;
sine[3173]=71;
sine[3174]=71;
sine[3175]=71;
sine[3176]=71;
sine[3177]=71;
sine[3178]=71;
sine[3179]=71;
sine[3180]=71;
sine[3181]=71;
sine[3182]=71;
sine[3183]=71;
sine[3184]=71;
sine[3185]=71;
sine[3186]=71;
sine[3187]=71;
sine[3188]=71;
sine[3189]=71;
sine[3190]=71;
sine[3191]=71;
sine[3192]=71;
sine[3193]=71;
sine[3194]=71;
sine[3195]=71;
sine[3196]=71;
sine[3197]=71;
sine[3198]=71;
sine[3199]=71;
sine[3200]=71;
sine[3201]=71;
sine[3202]=71;
sine[3203]=71;
sine[3204]=71;
sine[3205]=71;
sine[3206]=71;
sine[3207]=71;
sine[3208]=71;
sine[3209]=71;
sine[3210]=70;
sine[3211]=70;
sine[3212]=70;
sine[3213]=70;
sine[3214]=70;
sine[3215]=70;
sine[3216]=70;
sine[3217]=70;
sine[3218]=70;
sine[3219]=70;
sine[3220]=70;
sine[3221]=70;
sine[3222]=70;
sine[3223]=70;
sine[3224]=70;
sine[3225]=70;
sine[3226]=70;
sine[3227]=70;
sine[3228]=70;
sine[3229]=70;
sine[3230]=70;
sine[3231]=70;
sine[3232]=70;
sine[3233]=70;
sine[3234]=70;
sine[3235]=70;
sine[3236]=70;
sine[3237]=70;
sine[3238]=70;
sine[3239]=70;
sine[3240]=70;
sine[3241]=70;
sine[3242]=70;
sine[3243]=70;
sine[3244]=70;
sine[3245]=70;
sine[3246]=70;
sine[3247]=70;
sine[3248]=70;
sine[3249]=70;
sine[3250]=70;
sine[3251]=70;
sine[3252]=70;
sine[3253]=70;
sine[3254]=70;
sine[3255]=69;
sine[3256]=69;
sine[3257]=69;
sine[3258]=69;
sine[3259]=69;
sine[3260]=69;
sine[3261]=69;
sine[3262]=69;
sine[3263]=69;
sine[3264]=69;
sine[3265]=69;
sine[3266]=69;
sine[3267]=69;
sine[3268]=69;
sine[3269]=69;
sine[3270]=69;
sine[3271]=69;
sine[3272]=69;
sine[3273]=69;
sine[3274]=69;
sine[3275]=69;
sine[3276]=69;
sine[3277]=69;
sine[3278]=69;
sine[3279]=69;
sine[3280]=69;
sine[3281]=69;
sine[3282]=69;
sine[3283]=69;
sine[3284]=69;
sine[3285]=69;
sine[3286]=69;
sine[3287]=69;
sine[3288]=69;
sine[3289]=69;
sine[3290]=69;
sine[3291]=69;
sine[3292]=69;
sine[3293]=69;
sine[3294]=69;
sine[3295]=69;
sine[3296]=69;
sine[3297]=69;
sine[3298]=69;
sine[3299]=68;
sine[3300]=68;
sine[3301]=68;
sine[3302]=68;
sine[3303]=68;
sine[3304]=68;
sine[3305]=68;
sine[3306]=68;
sine[3307]=68;
sine[3308]=68;
sine[3309]=68;
sine[3310]=68;
sine[3311]=68;
sine[3312]=68;
sine[3313]=68;
sine[3314]=68;
sine[3315]=68;
sine[3316]=68;
sine[3317]=68;
sine[3318]=68;
sine[3319]=68;
sine[3320]=68;
sine[3321]=68;
sine[3322]=68;
sine[3323]=68;
sine[3324]=68;
sine[3325]=68;
sine[3326]=68;
sine[3327]=68;
sine[3328]=68;
sine[3329]=68;
sine[3330]=68;
sine[3331]=68;
sine[3332]=68;
sine[3333]=68;
sine[3334]=68;
sine[3335]=68;
sine[3336]=68;
sine[3337]=68;
sine[3338]=68;
sine[3339]=68;
sine[3340]=67;
sine[3341]=67;
sine[3342]=67;
sine[3343]=67;
sine[3344]=67;
sine[3345]=67;
sine[3346]=67;
sine[3347]=67;
sine[3348]=67;
sine[3349]=67;
sine[3350]=67;
sine[3351]=67;
sine[3352]=67;
sine[3353]=67;
sine[3354]=67;
sine[3355]=67;
sine[3356]=67;
sine[3357]=67;
sine[3358]=67;
sine[3359]=67;
sine[3360]=67;
sine[3361]=67;
sine[3362]=67;
sine[3363]=67;
sine[3364]=67;
sine[3365]=67;
sine[3366]=67;
sine[3367]=67;
sine[3368]=67;
sine[3369]=67;
sine[3370]=67;
sine[3371]=67;
sine[3372]=67;
sine[3373]=67;
sine[3374]=67;
sine[3375]=67;
sine[3376]=67;
sine[3377]=67;
sine[3378]=67;
sine[3379]=67;
sine[3380]=66;
sine[3381]=66;
sine[3382]=66;
sine[3383]=66;
sine[3384]=66;
sine[3385]=66;
sine[3386]=66;
sine[3387]=66;
sine[3388]=66;
sine[3389]=66;
sine[3390]=66;
sine[3391]=66;
sine[3392]=66;
sine[3393]=66;
sine[3394]=66;
sine[3395]=66;
sine[3396]=66;
sine[3397]=66;
sine[3398]=66;
sine[3399]=66;
sine[3400]=66;
sine[3401]=66;
sine[3402]=66;
sine[3403]=66;
sine[3404]=66;
sine[3405]=66;
sine[3406]=66;
sine[3407]=66;
sine[3408]=66;
sine[3409]=66;
sine[3410]=66;
sine[3411]=66;
sine[3412]=66;
sine[3413]=66;
sine[3414]=66;
sine[3415]=66;
sine[3416]=66;
sine[3417]=66;
sine[3418]=65;
sine[3419]=65;
sine[3420]=65;
sine[3421]=65;
sine[3422]=65;
sine[3423]=65;
sine[3424]=65;
sine[3425]=65;
sine[3426]=65;
sine[3427]=65;
sine[3428]=65;
sine[3429]=65;
sine[3430]=65;
sine[3431]=65;
sine[3432]=65;
sine[3433]=65;
sine[3434]=65;
sine[3435]=65;
sine[3436]=65;
sine[3437]=65;
sine[3438]=65;
sine[3439]=65;
sine[3440]=65;
sine[3441]=65;
sine[3442]=65;
sine[3443]=65;
sine[3444]=65;
sine[3445]=65;
sine[3446]=65;
sine[3447]=65;
sine[3448]=65;
sine[3449]=65;
sine[3450]=65;
sine[3451]=65;
sine[3452]=65;
sine[3453]=65;
sine[3454]=65;
sine[3455]=64;
sine[3456]=64;
sine[3457]=64;
sine[3458]=64;
sine[3459]=64;
sine[3460]=64;
sine[3461]=64;
sine[3462]=64;
sine[3463]=64;
sine[3464]=64;
sine[3465]=64;
sine[3466]=64;
sine[3467]=64;
sine[3468]=64;
sine[3469]=64;
sine[3470]=64;
sine[3471]=64;
sine[3472]=64;
sine[3473]=64;
sine[3474]=64;
sine[3475]=64;
sine[3476]=64;
sine[3477]=64;
sine[3478]=64;
sine[3479]=64;
sine[3480]=64;
sine[3481]=64;
sine[3482]=64;
sine[3483]=64;
sine[3484]=64;
sine[3485]=64;
sine[3486]=64;
sine[3487]=64;
sine[3488]=64;
sine[3489]=64;
sine[3490]=63;
sine[3491]=63;
sine[3492]=63;
sine[3493]=63;
sine[3494]=63;
sine[3495]=63;
sine[3496]=63;
sine[3497]=63;
sine[3498]=63;
sine[3499]=63;
sine[3500]=63;
sine[3501]=63;
sine[3502]=63;
sine[3503]=63;
sine[3504]=63;
sine[3505]=63;
sine[3506]=63;
sine[3507]=63;
sine[3508]=63;
sine[3509]=63;
sine[3510]=63;
sine[3511]=63;
sine[3512]=63;
sine[3513]=63;
sine[3514]=63;
sine[3515]=63;
sine[3516]=63;
sine[3517]=63;
sine[3518]=63;
sine[3519]=63;
sine[3520]=63;
sine[3521]=63;
sine[3522]=63;
sine[3523]=63;
sine[3524]=63;
sine[3525]=62;
sine[3526]=62;
sine[3527]=62;
sine[3528]=62;
sine[3529]=62;
sine[3530]=62;
sine[3531]=62;
sine[3532]=62;
sine[3533]=62;
sine[3534]=62;
sine[3535]=62;
sine[3536]=62;
sine[3537]=62;
sine[3538]=62;
sine[3539]=62;
sine[3540]=62;
sine[3541]=62;
sine[3542]=62;
sine[3543]=62;
sine[3544]=62;
sine[3545]=62;
sine[3546]=62;
sine[3547]=62;
sine[3548]=62;
sine[3549]=62;
sine[3550]=62;
sine[3551]=62;
sine[3552]=62;
sine[3553]=62;
sine[3554]=62;
sine[3555]=62;
sine[3556]=62;
sine[3557]=62;
sine[3558]=61;
sine[3559]=61;
sine[3560]=61;
sine[3561]=61;
sine[3562]=61;
sine[3563]=61;
sine[3564]=61;
sine[3565]=61;
sine[3566]=61;
sine[3567]=61;
sine[3568]=61;
sine[3569]=61;
sine[3570]=61;
sine[3571]=61;
sine[3572]=61;
sine[3573]=61;
sine[3574]=61;
sine[3575]=61;
sine[3576]=61;
sine[3577]=61;
sine[3578]=61;
sine[3579]=61;
sine[3580]=61;
sine[3581]=61;
sine[3582]=61;
sine[3583]=61;
sine[3584]=61;
sine[3585]=61;
sine[3586]=61;
sine[3587]=61;
sine[3588]=61;
sine[3589]=61;
sine[3590]=61;
sine[3591]=60;
sine[3592]=60;
sine[3593]=60;
sine[3594]=60;
sine[3595]=60;
sine[3596]=60;
sine[3597]=60;
sine[3598]=60;
sine[3599]=60;
sine[3600]=60;
sine[3601]=60;
sine[3602]=60;
sine[3603]=60;
sine[3604]=60;
sine[3605]=60;
sine[3606]=60;
sine[3607]=60;
sine[3608]=60;
sine[3609]=60;
sine[3610]=60;
sine[3611]=60;
sine[3612]=60;
sine[3613]=60;
sine[3614]=60;
sine[3615]=60;
sine[3616]=60;
sine[3617]=60;
sine[3618]=60;
sine[3619]=60;
sine[3620]=60;
sine[3621]=60;
sine[3622]=60;
sine[3623]=59;
sine[3624]=59;
sine[3625]=59;
sine[3626]=59;
sine[3627]=59;
sine[3628]=59;
sine[3629]=59;
sine[3630]=59;
sine[3631]=59;
sine[3632]=59;
sine[3633]=59;
sine[3634]=59;
sine[3635]=59;
sine[3636]=59;
sine[3637]=59;
sine[3638]=59;
sine[3639]=59;
sine[3640]=59;
sine[3641]=59;
sine[3642]=59;
sine[3643]=59;
sine[3644]=59;
sine[3645]=59;
sine[3646]=59;
sine[3647]=59;
sine[3648]=59;
sine[3649]=59;
sine[3650]=59;
sine[3651]=59;
sine[3652]=59;
sine[3653]=59;
sine[3654]=58;
sine[3655]=58;
sine[3656]=58;
sine[3657]=58;
sine[3658]=58;
sine[3659]=58;
sine[3660]=58;
sine[3661]=58;
sine[3662]=58;
sine[3663]=58;
sine[3664]=58;
sine[3665]=58;
sine[3666]=58;
sine[3667]=58;
sine[3668]=58;
sine[3669]=58;
sine[3670]=58;
sine[3671]=58;
sine[3672]=58;
sine[3673]=58;
sine[3674]=58;
sine[3675]=58;
sine[3676]=58;
sine[3677]=58;
sine[3678]=58;
sine[3679]=58;
sine[3680]=58;
sine[3681]=58;
sine[3682]=58;
sine[3683]=58;
sine[3684]=57;
sine[3685]=57;
sine[3686]=57;
sine[3687]=57;
sine[3688]=57;
sine[3689]=57;
sine[3690]=57;
sine[3691]=57;
sine[3692]=57;
sine[3693]=57;
sine[3694]=57;
sine[3695]=57;
sine[3696]=57;
sine[3697]=57;
sine[3698]=57;
sine[3699]=57;
sine[3700]=57;
sine[3701]=57;
sine[3702]=57;
sine[3703]=57;
sine[3704]=57;
sine[3705]=57;
sine[3706]=57;
sine[3707]=57;
sine[3708]=57;
sine[3709]=57;
sine[3710]=57;
sine[3711]=57;
sine[3712]=57;
sine[3713]=57;
sine[3714]=56;
sine[3715]=56;
sine[3716]=56;
sine[3717]=56;
sine[3718]=56;
sine[3719]=56;
sine[3720]=56;
sine[3721]=56;
sine[3722]=56;
sine[3723]=56;
sine[3724]=56;
sine[3725]=56;
sine[3726]=56;
sine[3727]=56;
sine[3728]=56;
sine[3729]=56;
sine[3730]=56;
sine[3731]=56;
sine[3732]=56;
sine[3733]=56;
sine[3734]=56;
sine[3735]=56;
sine[3736]=56;
sine[3737]=56;
sine[3738]=56;
sine[3739]=56;
sine[3740]=56;
sine[3741]=56;
sine[3742]=56;
sine[3743]=55;
sine[3744]=55;
sine[3745]=55;
sine[3746]=55;
sine[3747]=55;
sine[3748]=55;
sine[3749]=55;
sine[3750]=55;
sine[3751]=55;
sine[3752]=55;
sine[3753]=55;
sine[3754]=55;
sine[3755]=55;
sine[3756]=55;
sine[3757]=55;
sine[3758]=55;
sine[3759]=55;
sine[3760]=55;
sine[3761]=55;
sine[3762]=55;
sine[3763]=55;
sine[3764]=55;
sine[3765]=55;
sine[3766]=55;
sine[3767]=55;
sine[3768]=55;
sine[3769]=55;
sine[3770]=55;
sine[3771]=55;
sine[3772]=54;
sine[3773]=54;
sine[3774]=54;
sine[3775]=54;
sine[3776]=54;
sine[3777]=54;
sine[3778]=54;
sine[3779]=54;
sine[3780]=54;
sine[3781]=54;
sine[3782]=54;
sine[3783]=54;
sine[3784]=54;
sine[3785]=54;
sine[3786]=54;
sine[3787]=54;
sine[3788]=54;
sine[3789]=54;
sine[3790]=54;
sine[3791]=54;
sine[3792]=54;
sine[3793]=54;
sine[3794]=54;
sine[3795]=54;
sine[3796]=54;
sine[3797]=54;
sine[3798]=54;
sine[3799]=54;
sine[3800]=53;
sine[3801]=53;
sine[3802]=53;
sine[3803]=53;
sine[3804]=53;
sine[3805]=53;
sine[3806]=53;
sine[3807]=53;
sine[3808]=53;
sine[3809]=53;
sine[3810]=53;
sine[3811]=53;
sine[3812]=53;
sine[3813]=53;
sine[3814]=53;
sine[3815]=53;
sine[3816]=53;
sine[3817]=53;
sine[3818]=53;
sine[3819]=53;
sine[3820]=53;
sine[3821]=53;
sine[3822]=53;
sine[3823]=53;
sine[3824]=53;
sine[3825]=53;
sine[3826]=53;
sine[3827]=53;
sine[3828]=52;
sine[3829]=52;
sine[3830]=52;
sine[3831]=52;
sine[3832]=52;
sine[3833]=52;
sine[3834]=52;
sine[3835]=52;
sine[3836]=52;
sine[3837]=52;
sine[3838]=52;
sine[3839]=52;
sine[3840]=52;
sine[3841]=52;
sine[3842]=52;
sine[3843]=52;
sine[3844]=52;
sine[3845]=52;
sine[3846]=52;
sine[3847]=52;
sine[3848]=52;
sine[3849]=52;
sine[3850]=52;
sine[3851]=52;
sine[3852]=52;
sine[3853]=52;
sine[3854]=52;
sine[3855]=51;
sine[3856]=51;
sine[3857]=51;
sine[3858]=51;
sine[3859]=51;
sine[3860]=51;
sine[3861]=51;
sine[3862]=51;
sine[3863]=51;
sine[3864]=51;
sine[3865]=51;
sine[3866]=51;
sine[3867]=51;
sine[3868]=51;
sine[3869]=51;
sine[3870]=51;
sine[3871]=51;
sine[3872]=51;
sine[3873]=51;
sine[3874]=51;
sine[3875]=51;
sine[3876]=51;
sine[3877]=51;
sine[3878]=51;
sine[3879]=51;
sine[3880]=51;
sine[3881]=51;
sine[3882]=50;
sine[3883]=50;
sine[3884]=50;
sine[3885]=50;
sine[3886]=50;
sine[3887]=50;
sine[3888]=50;
sine[3889]=50;
sine[3890]=50;
sine[3891]=50;
sine[3892]=50;
sine[3893]=50;
sine[3894]=50;
sine[3895]=50;
sine[3896]=50;
sine[3897]=50;
sine[3898]=50;
sine[3899]=50;
sine[3900]=50;
sine[3901]=50;
sine[3902]=50;
sine[3903]=50;
sine[3904]=50;
sine[3905]=50;
sine[3906]=50;
sine[3907]=50;
sine[3908]=49;
sine[3909]=49;
sine[3910]=49;
sine[3911]=49;
sine[3912]=49;
sine[3913]=49;
sine[3914]=49;
sine[3915]=49;
sine[3916]=49;
sine[3917]=49;
sine[3918]=49;
sine[3919]=49;
sine[3920]=49;
sine[3921]=49;
sine[3922]=49;
sine[3923]=49;
sine[3924]=49;
sine[3925]=49;
sine[3926]=49;
sine[3927]=49;
sine[3928]=49;
sine[3929]=49;
sine[3930]=49;
sine[3931]=49;
sine[3932]=49;
sine[3933]=49;
sine[3934]=49;
sine[3935]=48;
sine[3936]=48;
sine[3937]=48;
sine[3938]=48;
sine[3939]=48;
sine[3940]=48;
sine[3941]=48;
sine[3942]=48;
sine[3943]=48;
sine[3944]=48;
sine[3945]=48;
sine[3946]=48;
sine[3947]=48;
sine[3948]=48;
sine[3949]=48;
sine[3950]=48;
sine[3951]=48;
sine[3952]=48;
sine[3953]=48;
sine[3954]=48;
sine[3955]=48;
sine[3956]=48;
sine[3957]=48;
sine[3958]=48;
sine[3959]=48;
sine[3960]=47;
sine[3961]=47;
sine[3962]=47;
sine[3963]=47;
sine[3964]=47;
sine[3965]=47;
sine[3966]=47;
sine[3967]=47;
sine[3968]=47;
sine[3969]=47;
sine[3970]=47;
sine[3971]=47;
sine[3972]=47;
sine[3973]=47;
sine[3974]=47;
sine[3975]=47;
sine[3976]=47;
sine[3977]=47;
sine[3978]=47;
sine[3979]=47;
sine[3980]=47;
sine[3981]=47;
sine[3982]=47;
sine[3983]=47;
sine[3984]=47;
sine[3985]=47;
sine[3986]=46;
sine[3987]=46;
sine[3988]=46;
sine[3989]=46;
sine[3990]=46;
sine[3991]=46;
sine[3992]=46;
sine[3993]=46;
sine[3994]=46;
sine[3995]=46;
sine[3996]=46;
sine[3997]=46;
sine[3998]=46;
sine[3999]=46;
sine[4000]=46;
sine[4001]=46;
sine[4002]=46;
sine[4003]=46;
sine[4004]=46;
sine[4005]=46;
sine[4006]=46;
sine[4007]=46;
sine[4008]=46;
sine[4009]=46;
sine[4010]=46;
sine[4011]=45;
sine[4012]=45;
sine[4013]=45;
sine[4014]=45;
sine[4015]=45;
sine[4016]=45;
sine[4017]=45;
sine[4018]=45;
sine[4019]=45;
sine[4020]=45;
sine[4021]=45;
sine[4022]=45;
sine[4023]=45;
sine[4024]=45;
sine[4025]=45;
sine[4026]=45;
sine[4027]=45;
sine[4028]=45;
sine[4029]=45;
sine[4030]=45;
sine[4031]=45;
sine[4032]=45;
sine[4033]=45;
sine[4034]=45;
sine[4035]=45;
sine[4036]=44;
sine[4037]=44;
sine[4038]=44;
sine[4039]=44;
sine[4040]=44;
sine[4041]=44;
sine[4042]=44;
sine[4043]=44;
sine[4044]=44;
sine[4045]=44;
sine[4046]=44;
sine[4047]=44;
sine[4048]=44;
sine[4049]=44;
sine[4050]=44;
sine[4051]=44;
sine[4052]=44;
sine[4053]=44;
sine[4054]=44;
sine[4055]=44;
sine[4056]=44;
sine[4057]=44;
sine[4058]=44;
sine[4059]=44;
sine[4060]=44;
sine[4061]=43;
sine[4062]=43;
sine[4063]=43;
sine[4064]=43;
sine[4065]=43;
sine[4066]=43;
sine[4067]=43;
sine[4068]=43;
sine[4069]=43;
sine[4070]=43;
sine[4071]=43;
sine[4072]=43;
sine[4073]=43;
sine[4074]=43;
sine[4075]=43;
sine[4076]=43;
sine[4077]=43;
sine[4078]=43;
sine[4079]=43;
sine[4080]=43;
sine[4081]=43;
sine[4082]=43;
sine[4083]=43;
sine[4084]=43;
sine[4085]=42;
sine[4086]=42;
sine[4087]=42;
sine[4088]=42;
sine[4089]=42;
sine[4090]=42;
sine[4091]=42;
sine[4092]=42;
sine[4093]=42;
sine[4094]=42;
sine[4095]=42;
sine[4096]=42;
sine[4097]=42;
sine[4098]=42;
sine[4099]=42;
sine[4100]=42;
sine[4101]=42;
sine[4102]=42;
sine[4103]=42;
sine[4104]=42;
sine[4105]=42;
sine[4106]=42;
sine[4107]=42;
sine[4108]=42;
sine[4109]=41;
sine[4110]=41;
sine[4111]=41;
sine[4112]=41;
sine[4113]=41;
sine[4114]=41;
sine[4115]=41;
sine[4116]=41;
sine[4117]=41;
sine[4118]=41;
sine[4119]=41;
sine[4120]=41;
sine[4121]=41;
sine[4122]=41;
sine[4123]=41;
sine[4124]=41;
sine[4125]=41;
sine[4126]=41;
sine[4127]=41;
sine[4128]=41;
sine[4129]=41;
sine[4130]=41;
sine[4131]=41;
sine[4132]=41;
sine[4133]=40;
sine[4134]=40;
sine[4135]=40;
sine[4136]=40;
sine[4137]=40;
sine[4138]=40;
sine[4139]=40;
sine[4140]=40;
sine[4141]=40;
sine[4142]=40;
sine[4143]=40;
sine[4144]=40;
sine[4145]=40;
sine[4146]=40;
sine[4147]=40;
sine[4148]=40;
sine[4149]=40;
sine[4150]=40;
sine[4151]=40;
sine[4152]=40;
sine[4153]=40;
sine[4154]=40;
sine[4155]=40;
sine[4156]=40;
sine[4157]=39;
sine[4158]=39;
sine[4159]=39;
sine[4160]=39;
sine[4161]=39;
sine[4162]=39;
sine[4163]=39;
sine[4164]=39;
sine[4165]=39;
sine[4166]=39;
sine[4167]=39;
sine[4168]=39;
sine[4169]=39;
sine[4170]=39;
sine[4171]=39;
sine[4172]=39;
sine[4173]=39;
sine[4174]=39;
sine[4175]=39;
sine[4176]=39;
sine[4177]=39;
sine[4178]=39;
sine[4179]=39;
sine[4180]=38;
sine[4181]=38;
sine[4182]=38;
sine[4183]=38;
sine[4184]=38;
sine[4185]=38;
sine[4186]=38;
sine[4187]=38;
sine[4188]=38;
sine[4189]=38;
sine[4190]=38;
sine[4191]=38;
sine[4192]=38;
sine[4193]=38;
sine[4194]=38;
sine[4195]=38;
sine[4196]=38;
sine[4197]=38;
sine[4198]=38;
sine[4199]=38;
sine[4200]=38;
sine[4201]=38;
sine[4202]=38;
sine[4203]=38;
sine[4204]=37;
sine[4205]=37;
sine[4206]=37;
sine[4207]=37;
sine[4208]=37;
sine[4209]=37;
sine[4210]=37;
sine[4211]=37;
sine[4212]=37;
sine[4213]=37;
sine[4214]=37;
sine[4215]=37;
sine[4216]=37;
sine[4217]=37;
sine[4218]=37;
sine[4219]=37;
sine[4220]=37;
sine[4221]=37;
sine[4222]=37;
sine[4223]=37;
sine[4224]=37;
sine[4225]=37;
sine[4226]=37;
sine[4227]=36;
sine[4228]=36;
sine[4229]=36;
sine[4230]=36;
sine[4231]=36;
sine[4232]=36;
sine[4233]=36;
sine[4234]=36;
sine[4235]=36;
sine[4236]=36;
sine[4237]=36;
sine[4238]=36;
sine[4239]=36;
sine[4240]=36;
sine[4241]=36;
sine[4242]=36;
sine[4243]=36;
sine[4244]=36;
sine[4245]=36;
sine[4246]=36;
sine[4247]=36;
sine[4248]=36;
sine[4249]=36;
sine[4250]=35;
sine[4251]=35;
sine[4252]=35;
sine[4253]=35;
sine[4254]=35;
sine[4255]=35;
sine[4256]=35;
sine[4257]=35;
sine[4258]=35;
sine[4259]=35;
sine[4260]=35;
sine[4261]=35;
sine[4262]=35;
sine[4263]=35;
sine[4264]=35;
sine[4265]=35;
sine[4266]=35;
sine[4267]=35;
sine[4268]=35;
sine[4269]=35;
sine[4270]=35;
sine[4271]=35;
sine[4272]=35;
sine[4273]=34;
sine[4274]=34;
sine[4275]=34;
sine[4276]=34;
sine[4277]=34;
sine[4278]=34;
sine[4279]=34;
sine[4280]=34;
sine[4281]=34;
sine[4282]=34;
sine[4283]=34;
sine[4284]=34;
sine[4285]=34;
sine[4286]=34;
sine[4287]=34;
sine[4288]=34;
sine[4289]=34;
sine[4290]=34;
sine[4291]=34;
sine[4292]=34;
sine[4293]=34;
sine[4294]=34;
sine[4295]=33;
sine[4296]=33;
sine[4297]=33;
sine[4298]=33;
sine[4299]=33;
sine[4300]=33;
sine[4301]=33;
sine[4302]=33;
sine[4303]=33;
sine[4304]=33;
sine[4305]=33;
sine[4306]=33;
sine[4307]=33;
sine[4308]=33;
sine[4309]=33;
sine[4310]=33;
sine[4311]=33;
sine[4312]=33;
sine[4313]=33;
sine[4314]=33;
sine[4315]=33;
sine[4316]=33;
sine[4317]=33;
sine[4318]=32;
sine[4319]=32;
sine[4320]=32;
sine[4321]=32;
sine[4322]=32;
sine[4323]=32;
sine[4324]=32;
sine[4325]=32;
sine[4326]=32;
sine[4327]=32;
sine[4328]=32;
sine[4329]=32;
sine[4330]=32;
sine[4331]=32;
sine[4332]=32;
sine[4333]=32;
sine[4334]=32;
sine[4335]=32;
sine[4336]=32;
sine[4337]=32;
sine[4338]=32;
sine[4339]=32;
sine[4340]=31;
sine[4341]=31;
sine[4342]=31;
sine[4343]=31;
sine[4344]=31;
sine[4345]=31;
sine[4346]=31;
sine[4347]=31;
sine[4348]=31;
sine[4349]=31;
sine[4350]=31;
sine[4351]=31;
sine[4352]=31;
sine[4353]=31;
sine[4354]=31;
sine[4355]=31;
sine[4356]=31;
sine[4357]=31;
sine[4358]=31;
sine[4359]=31;
sine[4360]=31;
sine[4361]=31;
sine[4362]=30;
sine[4363]=30;
sine[4364]=30;
sine[4365]=30;
sine[4366]=30;
sine[4367]=30;
sine[4368]=30;
sine[4369]=30;
sine[4370]=30;
sine[4371]=30;
sine[4372]=30;
sine[4373]=30;
sine[4374]=30;
sine[4375]=30;
sine[4376]=30;
sine[4377]=30;
sine[4378]=30;
sine[4379]=30;
sine[4380]=30;
sine[4381]=30;
sine[4382]=30;
sine[4383]=30;
sine[4384]=29;
sine[4385]=29;
sine[4386]=29;
sine[4387]=29;
sine[4388]=29;
sine[4389]=29;
sine[4390]=29;
sine[4391]=29;
sine[4392]=29;
sine[4393]=29;
sine[4394]=29;
sine[4395]=29;
sine[4396]=29;
sine[4397]=29;
sine[4398]=29;
sine[4399]=29;
sine[4400]=29;
sine[4401]=29;
sine[4402]=29;
sine[4403]=29;
sine[4404]=29;
sine[4405]=29;
sine[4406]=28;
sine[4407]=28;
sine[4408]=28;
sine[4409]=28;
sine[4410]=28;
sine[4411]=28;
sine[4412]=28;
sine[4413]=28;
sine[4414]=28;
sine[4415]=28;
sine[4416]=28;
sine[4417]=28;
sine[4418]=28;
sine[4419]=28;
sine[4420]=28;
sine[4421]=28;
sine[4422]=28;
sine[4423]=28;
sine[4424]=28;
sine[4425]=28;
sine[4426]=28;
sine[4427]=28;
sine[4428]=27;
sine[4429]=27;
sine[4430]=27;
sine[4431]=27;
sine[4432]=27;
sine[4433]=27;
sine[4434]=27;
sine[4435]=27;
sine[4436]=27;
sine[4437]=27;
sine[4438]=27;
sine[4439]=27;
sine[4440]=27;
sine[4441]=27;
sine[4442]=27;
sine[4443]=27;
sine[4444]=27;
sine[4445]=27;
sine[4446]=27;
sine[4447]=27;
sine[4448]=27;
sine[4449]=27;
sine[4450]=26;
sine[4451]=26;
sine[4452]=26;
sine[4453]=26;
sine[4454]=26;
sine[4455]=26;
sine[4456]=26;
sine[4457]=26;
sine[4458]=26;
sine[4459]=26;
sine[4460]=26;
sine[4461]=26;
sine[4462]=26;
sine[4463]=26;
sine[4464]=26;
sine[4465]=26;
sine[4466]=26;
sine[4467]=26;
sine[4468]=26;
sine[4469]=26;
sine[4470]=26;
sine[4471]=25;
sine[4472]=25;
sine[4473]=25;
sine[4474]=25;
sine[4475]=25;
sine[4476]=25;
sine[4477]=25;
sine[4478]=25;
sine[4479]=25;
sine[4480]=25;
sine[4481]=25;
sine[4482]=25;
sine[4483]=25;
sine[4484]=25;
sine[4485]=25;
sine[4486]=25;
sine[4487]=25;
sine[4488]=25;
sine[4489]=25;
sine[4490]=25;
sine[4491]=25;
sine[4492]=25;
sine[4493]=24;
sine[4494]=24;
sine[4495]=24;
sine[4496]=24;
sine[4497]=24;
sine[4498]=24;
sine[4499]=24;
sine[4500]=24;
sine[4501]=24;
sine[4502]=24;
sine[4503]=24;
sine[4504]=24;
sine[4505]=24;
sine[4506]=24;
sine[4507]=24;
sine[4508]=24;
sine[4509]=24;
sine[4510]=24;
sine[4511]=24;
sine[4512]=24;
sine[4513]=24;
sine[4514]=23;
sine[4515]=23;
sine[4516]=23;
sine[4517]=23;
sine[4518]=23;
sine[4519]=23;
sine[4520]=23;
sine[4521]=23;
sine[4522]=23;
sine[4523]=23;
sine[4524]=23;
sine[4525]=23;
sine[4526]=23;
sine[4527]=23;
sine[4528]=23;
sine[4529]=23;
sine[4530]=23;
sine[4531]=23;
sine[4532]=23;
sine[4533]=23;
sine[4534]=23;
sine[4535]=23;
sine[4536]=22;
sine[4537]=22;
sine[4538]=22;
sine[4539]=22;
sine[4540]=22;
sine[4541]=22;
sine[4542]=22;
sine[4543]=22;
sine[4544]=22;
sine[4545]=22;
sine[4546]=22;
sine[4547]=22;
sine[4548]=22;
sine[4549]=22;
sine[4550]=22;
sine[4551]=22;
sine[4552]=22;
sine[4553]=22;
sine[4554]=22;
sine[4555]=22;
sine[4556]=22;
sine[4557]=21;
sine[4558]=21;
sine[4559]=21;
sine[4560]=21;
sine[4561]=21;
sine[4562]=21;
sine[4563]=21;
sine[4564]=21;
sine[4565]=21;
sine[4566]=21;
sine[4567]=21;
sine[4568]=21;
sine[4569]=21;
sine[4570]=21;
sine[4571]=21;
sine[4572]=21;
sine[4573]=21;
sine[4574]=21;
sine[4575]=21;
sine[4576]=21;
sine[4577]=21;
sine[4578]=20;
sine[4579]=20;
sine[4580]=20;
sine[4581]=20;
sine[4582]=20;
sine[4583]=20;
sine[4584]=20;
sine[4585]=20;
sine[4586]=20;
sine[4587]=20;
sine[4588]=20;
sine[4589]=20;
sine[4590]=20;
sine[4591]=20;
sine[4592]=20;
sine[4593]=20;
sine[4594]=20;
sine[4595]=20;
sine[4596]=20;
sine[4597]=20;
sine[4598]=20;
sine[4599]=19;
sine[4600]=19;
sine[4601]=19;
sine[4602]=19;
sine[4603]=19;
sine[4604]=19;
sine[4605]=19;
sine[4606]=19;
sine[4607]=19;
sine[4608]=19;
sine[4609]=19;
sine[4610]=19;
sine[4611]=19;
sine[4612]=19;
sine[4613]=19;
sine[4614]=19;
sine[4615]=19;
sine[4616]=19;
sine[4617]=19;
sine[4618]=19;
sine[4619]=19;
sine[4620]=18;
sine[4621]=18;
sine[4622]=18;
sine[4623]=18;
sine[4624]=18;
sine[4625]=18;
sine[4626]=18;
sine[4627]=18;
sine[4628]=18;
sine[4629]=18;
sine[4630]=18;
sine[4631]=18;
sine[4632]=18;
sine[4633]=18;
sine[4634]=18;
sine[4635]=18;
sine[4636]=18;
sine[4637]=18;
sine[4638]=18;
sine[4639]=18;
sine[4640]=18;
sine[4641]=17;
sine[4642]=17;
sine[4643]=17;
sine[4644]=17;
sine[4645]=17;
sine[4646]=17;
sine[4647]=17;
sine[4648]=17;
sine[4649]=17;
sine[4650]=17;
sine[4651]=17;
sine[4652]=17;
sine[4653]=17;
sine[4654]=17;
sine[4655]=17;
sine[4656]=17;
sine[4657]=17;
sine[4658]=17;
sine[4659]=17;
sine[4660]=17;
sine[4661]=17;
sine[4662]=16;
sine[4663]=16;
sine[4664]=16;
sine[4665]=16;
sine[4666]=16;
sine[4667]=16;
sine[4668]=16;
sine[4669]=16;
sine[4670]=16;
sine[4671]=16;
sine[4672]=16;
sine[4673]=16;
sine[4674]=16;
sine[4675]=16;
sine[4676]=16;
sine[4677]=16;
sine[4678]=16;
sine[4679]=16;
sine[4680]=16;
sine[4681]=16;
sine[4682]=16;
sine[4683]=15;
sine[4684]=15;
sine[4685]=15;
sine[4686]=15;
sine[4687]=15;
sine[4688]=15;
sine[4689]=15;
sine[4690]=15;
sine[4691]=15;
sine[4692]=15;
sine[4693]=15;
sine[4694]=15;
sine[4695]=15;
sine[4696]=15;
sine[4697]=15;
sine[4698]=15;
sine[4699]=15;
sine[4700]=15;
sine[4701]=15;
sine[4702]=15;
sine[4703]=14;
sine[4704]=14;
sine[4705]=14;
sine[4706]=14;
sine[4707]=14;
sine[4708]=14;
sine[4709]=14;
sine[4710]=14;
sine[4711]=14;
sine[4712]=14;
sine[4713]=14;
sine[4714]=14;
sine[4715]=14;
sine[4716]=14;
sine[4717]=14;
sine[4718]=14;
sine[4719]=14;
sine[4720]=14;
sine[4721]=14;
sine[4722]=14;
sine[4723]=14;
sine[4724]=13;
sine[4725]=13;
sine[4726]=13;
sine[4727]=13;
sine[4728]=13;
sine[4729]=13;
sine[4730]=13;
sine[4731]=13;
sine[4732]=13;
sine[4733]=13;
sine[4734]=13;
sine[4735]=13;
sine[4736]=13;
sine[4737]=13;
sine[4738]=13;
sine[4739]=13;
sine[4740]=13;
sine[4741]=13;
sine[4742]=13;
sine[4743]=13;
sine[4744]=13;
sine[4745]=12;
sine[4746]=12;
sine[4747]=12;
sine[4748]=12;
sine[4749]=12;
sine[4750]=12;
sine[4751]=12;
sine[4752]=12;
sine[4753]=12;
sine[4754]=12;
sine[4755]=12;
sine[4756]=12;
sine[4757]=12;
sine[4758]=12;
sine[4759]=12;
sine[4760]=12;
sine[4761]=12;
sine[4762]=12;
sine[4763]=12;
sine[4764]=12;
sine[4765]=11;
sine[4766]=11;
sine[4767]=11;
sine[4768]=11;
sine[4769]=11;
sine[4770]=11;
sine[4771]=11;
sine[4772]=11;
sine[4773]=11;
sine[4774]=11;
sine[4775]=11;
sine[4776]=11;
sine[4777]=11;
sine[4778]=11;
sine[4779]=11;
sine[4780]=11;
sine[4781]=11;
sine[4782]=11;
sine[4783]=11;
sine[4784]=11;
sine[4785]=11;
sine[4786]=10;
sine[4787]=10;
sine[4788]=10;
sine[4789]=10;
sine[4790]=10;
sine[4791]=10;
sine[4792]=10;
sine[4793]=10;
sine[4794]=10;
sine[4795]=10;
sine[4796]=10;
sine[4797]=10;
sine[4798]=10;
sine[4799]=10;
sine[4800]=10;
sine[4801]=10;
sine[4802]=10;
sine[4803]=10;
sine[4804]=10;
sine[4805]=10;
sine[4806]=9;
sine[4807]=9;
sine[4808]=9;
sine[4809]=9;
sine[4810]=9;
sine[4811]=9;
sine[4812]=9;
sine[4813]=9;
sine[4814]=9;
sine[4815]=9;
sine[4816]=9;
sine[4817]=9;
sine[4818]=9;
sine[4819]=9;
sine[4820]=9;
sine[4821]=9;
sine[4822]=9;
sine[4823]=9;
sine[4824]=9;
sine[4825]=9;
sine[4826]=9;
sine[4827]=8;
sine[4828]=8;
sine[4829]=8;
sine[4830]=8;
sine[4831]=8;
sine[4832]=8;
sine[4833]=8;
sine[4834]=8;
sine[4835]=8;
sine[4836]=8;
sine[4837]=8;
sine[4838]=8;
sine[4839]=8;
sine[4840]=8;
sine[4841]=8;
sine[4842]=8;
sine[4843]=8;
sine[4844]=8;
sine[4845]=8;
sine[4846]=8;
sine[4847]=7;
sine[4848]=7;
sine[4849]=7;
sine[4850]=7;
sine[4851]=7;
sine[4852]=7;
sine[4853]=7;
sine[4854]=7;
sine[4855]=7;
sine[4856]=7;
sine[4857]=7;
sine[4858]=7;
sine[4859]=7;
sine[4860]=7;
sine[4861]=7;
sine[4862]=7;
sine[4863]=7;
sine[4864]=7;
sine[4865]=7;
sine[4866]=7;
sine[4867]=7;
sine[4868]=6;
sine[4869]=6;
sine[4870]=6;
sine[4871]=6;
sine[4872]=6;
sine[4873]=6;
sine[4874]=6;
sine[4875]=6;
sine[4876]=6;
sine[4877]=6;
sine[4878]=6;
sine[4879]=6;
sine[4880]=6;
sine[4881]=6;
sine[4882]=6;
sine[4883]=6;
sine[4884]=6;
sine[4885]=6;
sine[4886]=6;
sine[4887]=6;
sine[4888]=5;
sine[4889]=5;
sine[4890]=5;
sine[4891]=5;
sine[4892]=5;
sine[4893]=5;
sine[4894]=5;
sine[4895]=5;
sine[4896]=5;
sine[4897]=5;
sine[4898]=5;
sine[4899]=5;
sine[4900]=5;
sine[4901]=5;
sine[4902]=5;
sine[4903]=5;
sine[4904]=5;
sine[4905]=5;
sine[4906]=5;
sine[4907]=5;
sine[4908]=5;
sine[4909]=4;
sine[4910]=4;
sine[4911]=4;
sine[4912]=4;
sine[4913]=4;
sine[4914]=4;
sine[4915]=4;
sine[4916]=4;
sine[4917]=4;
sine[4918]=4;
sine[4919]=4;
sine[4920]=4;
sine[4921]=4;
sine[4922]=4;
sine[4923]=4;
sine[4924]=4;
sine[4925]=4;
sine[4926]=4;
sine[4927]=4;
sine[4928]=4;
sine[4929]=3;
sine[4930]=3;
sine[4931]=3;
sine[4932]=3;
sine[4933]=3;
sine[4934]=3;
sine[4935]=3;
sine[4936]=3;
sine[4937]=3;
sine[4938]=3;
sine[4939]=3;
sine[4940]=3;
sine[4941]=3;
sine[4942]=3;
sine[4943]=3;
sine[4944]=3;
sine[4945]=3;
sine[4946]=3;
sine[4947]=3;
sine[4948]=3;
sine[4949]=3;
sine[4950]=2;
sine[4951]=2;
sine[4952]=2;
sine[4953]=2;
sine[4954]=2;
sine[4955]=2;
sine[4956]=2;
sine[4957]=2;
sine[4958]=2;
sine[4959]=2;
sine[4960]=2;
sine[4961]=2;
sine[4962]=2;
sine[4963]=2;
sine[4964]=2;
sine[4965]=2;
sine[4966]=2;
sine[4967]=2;
sine[4968]=2;
sine[4969]=2;
sine[4970]=1;
sine[4971]=1;
sine[4972]=1;
sine[4973]=1;
sine[4974]=1;
sine[4975]=1;
sine[4976]=1;
sine[4977]=1;
sine[4978]=1;
sine[4979]=1;
sine[4980]=1;
sine[4981]=1;
sine[4982]=1;
sine[4983]=1;
sine[4984]=1;
sine[4985]=1;
sine[4986]=1;
sine[4987]=1;
sine[4988]=1;
sine[4989]=1;
sine[4990]=0;
sine[4991]=0;
sine[4992]=0;
sine[4993]=0;
sine[4994]=0;
sine[4995]=0;
sine[4996]=0;
sine[4997]=0;
sine[4998]=0;
sine[4999]=0;
sine[5000]=0;
sine[5001]=0;
sine[5002]=0;
sine[5003]=0;
sine[5004]=0;
sine[5005]=0;
sine[5006]=0;
sine[5007]=0;
sine[5008]=0;
sine[5009]=0;
sine[5010]=0;
sine[5011]=-1;
sine[5012]=-1;
sine[5013]=-1;
sine[5014]=-1;
sine[5015]=-1;
sine[5016]=-1;
sine[5017]=-1;
sine[5018]=-1;
sine[5019]=-1;
sine[5020]=-1;
sine[5021]=-1;
sine[5022]=-1;
sine[5023]=-1;
sine[5024]=-1;
sine[5025]=-1;
sine[5026]=-1;
sine[5027]=-1;
sine[5028]=-1;
sine[5029]=-1;
sine[5030]=-1;
sine[5031]=-2;
sine[5032]=-2;
sine[5033]=-2;
sine[5034]=-2;
sine[5035]=-2;
sine[5036]=-2;
sine[5037]=-2;
sine[5038]=-2;
sine[5039]=-2;
sine[5040]=-2;
sine[5041]=-2;
sine[5042]=-2;
sine[5043]=-2;
sine[5044]=-2;
sine[5045]=-2;
sine[5046]=-2;
sine[5047]=-2;
sine[5048]=-2;
sine[5049]=-2;
sine[5050]=-2;
sine[5051]=-3;
sine[5052]=-3;
sine[5053]=-3;
sine[5054]=-3;
sine[5055]=-3;
sine[5056]=-3;
sine[5057]=-3;
sine[5058]=-3;
sine[5059]=-3;
sine[5060]=-3;
sine[5061]=-3;
sine[5062]=-3;
sine[5063]=-3;
sine[5064]=-3;
sine[5065]=-3;
sine[5066]=-3;
sine[5067]=-3;
sine[5068]=-3;
sine[5069]=-3;
sine[5070]=-3;
sine[5071]=-3;
sine[5072]=-4;
sine[5073]=-4;
sine[5074]=-4;
sine[5075]=-4;
sine[5076]=-4;
sine[5077]=-4;
sine[5078]=-4;
sine[5079]=-4;
sine[5080]=-4;
sine[5081]=-4;
sine[5082]=-4;
sine[5083]=-4;
sine[5084]=-4;
sine[5085]=-4;
sine[5086]=-4;
sine[5087]=-4;
sine[5088]=-4;
sine[5089]=-4;
sine[5090]=-4;
sine[5091]=-4;
sine[5092]=-5;
sine[5093]=-5;
sine[5094]=-5;
sine[5095]=-5;
sine[5096]=-5;
sine[5097]=-5;
sine[5098]=-5;
sine[5099]=-5;
sine[5100]=-5;
sine[5101]=-5;
sine[5102]=-5;
sine[5103]=-5;
sine[5104]=-5;
sine[5105]=-5;
sine[5106]=-5;
sine[5107]=-5;
sine[5108]=-5;
sine[5109]=-5;
sine[5110]=-5;
sine[5111]=-5;
sine[5112]=-5;
sine[5113]=-6;
sine[5114]=-6;
sine[5115]=-6;
sine[5116]=-6;
sine[5117]=-6;
sine[5118]=-6;
sine[5119]=-6;
sine[5120]=-6;
sine[5121]=-6;
sine[5122]=-6;
sine[5123]=-6;
sine[5124]=-6;
sine[5125]=-6;
sine[5126]=-6;
sine[5127]=-6;
sine[5128]=-6;
sine[5129]=-6;
sine[5130]=-6;
sine[5131]=-6;
sine[5132]=-6;
sine[5133]=-7;
sine[5134]=-7;
sine[5135]=-7;
sine[5136]=-7;
sine[5137]=-7;
sine[5138]=-7;
sine[5139]=-7;
sine[5140]=-7;
sine[5141]=-7;
sine[5142]=-7;
sine[5143]=-7;
sine[5144]=-7;
sine[5145]=-7;
sine[5146]=-7;
sine[5147]=-7;
sine[5148]=-7;
sine[5149]=-7;
sine[5150]=-7;
sine[5151]=-7;
sine[5152]=-7;
sine[5153]=-7;
sine[5154]=-8;
sine[5155]=-8;
sine[5156]=-8;
sine[5157]=-8;
sine[5158]=-8;
sine[5159]=-8;
sine[5160]=-8;
sine[5161]=-8;
sine[5162]=-8;
sine[5163]=-8;
sine[5164]=-8;
sine[5165]=-8;
sine[5166]=-8;
sine[5167]=-8;
sine[5168]=-8;
sine[5169]=-8;
sine[5170]=-8;
sine[5171]=-8;
sine[5172]=-8;
sine[5173]=-8;
sine[5174]=-9;
sine[5175]=-9;
sine[5176]=-9;
sine[5177]=-9;
sine[5178]=-9;
sine[5179]=-9;
sine[5180]=-9;
sine[5181]=-9;
sine[5182]=-9;
sine[5183]=-9;
sine[5184]=-9;
sine[5185]=-9;
sine[5186]=-9;
sine[5187]=-9;
sine[5188]=-9;
sine[5189]=-9;
sine[5190]=-9;
sine[5191]=-9;
sine[5192]=-9;
sine[5193]=-9;
sine[5194]=-9;
sine[5195]=-10;
sine[5196]=-10;
sine[5197]=-10;
sine[5198]=-10;
sine[5199]=-10;
sine[5200]=-10;
sine[5201]=-10;
sine[5202]=-10;
sine[5203]=-10;
sine[5204]=-10;
sine[5205]=-10;
sine[5206]=-10;
sine[5207]=-10;
sine[5208]=-10;
sine[5209]=-10;
sine[5210]=-10;
sine[5211]=-10;
sine[5212]=-10;
sine[5213]=-10;
sine[5214]=-10;
sine[5215]=-11;
sine[5216]=-11;
sine[5217]=-11;
sine[5218]=-11;
sine[5219]=-11;
sine[5220]=-11;
sine[5221]=-11;
sine[5222]=-11;
sine[5223]=-11;
sine[5224]=-11;
sine[5225]=-11;
sine[5226]=-11;
sine[5227]=-11;
sine[5228]=-11;
sine[5229]=-11;
sine[5230]=-11;
sine[5231]=-11;
sine[5232]=-11;
sine[5233]=-11;
sine[5234]=-11;
sine[5235]=-11;
sine[5236]=-12;
sine[5237]=-12;
sine[5238]=-12;
sine[5239]=-12;
sine[5240]=-12;
sine[5241]=-12;
sine[5242]=-12;
sine[5243]=-12;
sine[5244]=-12;
sine[5245]=-12;
sine[5246]=-12;
sine[5247]=-12;
sine[5248]=-12;
sine[5249]=-12;
sine[5250]=-12;
sine[5251]=-12;
sine[5252]=-12;
sine[5253]=-12;
sine[5254]=-12;
sine[5255]=-12;
sine[5256]=-13;
sine[5257]=-13;
sine[5258]=-13;
sine[5259]=-13;
sine[5260]=-13;
sine[5261]=-13;
sine[5262]=-13;
sine[5263]=-13;
sine[5264]=-13;
sine[5265]=-13;
sine[5266]=-13;
sine[5267]=-13;
sine[5268]=-13;
sine[5269]=-13;
sine[5270]=-13;
sine[5271]=-13;
sine[5272]=-13;
sine[5273]=-13;
sine[5274]=-13;
sine[5275]=-13;
sine[5276]=-13;
sine[5277]=-14;
sine[5278]=-14;
sine[5279]=-14;
sine[5280]=-14;
sine[5281]=-14;
sine[5282]=-14;
sine[5283]=-14;
sine[5284]=-14;
sine[5285]=-14;
sine[5286]=-14;
sine[5287]=-14;
sine[5288]=-14;
sine[5289]=-14;
sine[5290]=-14;
sine[5291]=-14;
sine[5292]=-14;
sine[5293]=-14;
sine[5294]=-14;
sine[5295]=-14;
sine[5296]=-14;
sine[5297]=-14;
sine[5298]=-15;
sine[5299]=-15;
sine[5300]=-15;
sine[5301]=-15;
sine[5302]=-15;
sine[5303]=-15;
sine[5304]=-15;
sine[5305]=-15;
sine[5306]=-15;
sine[5307]=-15;
sine[5308]=-15;
sine[5309]=-15;
sine[5310]=-15;
sine[5311]=-15;
sine[5312]=-15;
sine[5313]=-15;
sine[5314]=-15;
sine[5315]=-15;
sine[5316]=-15;
sine[5317]=-15;
sine[5318]=-16;
sine[5319]=-16;
sine[5320]=-16;
sine[5321]=-16;
sine[5322]=-16;
sine[5323]=-16;
sine[5324]=-16;
sine[5325]=-16;
sine[5326]=-16;
sine[5327]=-16;
sine[5328]=-16;
sine[5329]=-16;
sine[5330]=-16;
sine[5331]=-16;
sine[5332]=-16;
sine[5333]=-16;
sine[5334]=-16;
sine[5335]=-16;
sine[5336]=-16;
sine[5337]=-16;
sine[5338]=-16;
sine[5339]=-17;
sine[5340]=-17;
sine[5341]=-17;
sine[5342]=-17;
sine[5343]=-17;
sine[5344]=-17;
sine[5345]=-17;
sine[5346]=-17;
sine[5347]=-17;
sine[5348]=-17;
sine[5349]=-17;
sine[5350]=-17;
sine[5351]=-17;
sine[5352]=-17;
sine[5353]=-17;
sine[5354]=-17;
sine[5355]=-17;
sine[5356]=-17;
sine[5357]=-17;
sine[5358]=-17;
sine[5359]=-17;
sine[5360]=-18;
sine[5361]=-18;
sine[5362]=-18;
sine[5363]=-18;
sine[5364]=-18;
sine[5365]=-18;
sine[5366]=-18;
sine[5367]=-18;
sine[5368]=-18;
sine[5369]=-18;
sine[5370]=-18;
sine[5371]=-18;
sine[5372]=-18;
sine[5373]=-18;
sine[5374]=-18;
sine[5375]=-18;
sine[5376]=-18;
sine[5377]=-18;
sine[5378]=-18;
sine[5379]=-18;
sine[5380]=-18;
sine[5381]=-19;
sine[5382]=-19;
sine[5383]=-19;
sine[5384]=-19;
sine[5385]=-19;
sine[5386]=-19;
sine[5387]=-19;
sine[5388]=-19;
sine[5389]=-19;
sine[5390]=-19;
sine[5391]=-19;
sine[5392]=-19;
sine[5393]=-19;
sine[5394]=-19;
sine[5395]=-19;
sine[5396]=-19;
sine[5397]=-19;
sine[5398]=-19;
sine[5399]=-19;
sine[5400]=-19;
sine[5401]=-19;
sine[5402]=-20;
sine[5403]=-20;
sine[5404]=-20;
sine[5405]=-20;
sine[5406]=-20;
sine[5407]=-20;
sine[5408]=-20;
sine[5409]=-20;
sine[5410]=-20;
sine[5411]=-20;
sine[5412]=-20;
sine[5413]=-20;
sine[5414]=-20;
sine[5415]=-20;
sine[5416]=-20;
sine[5417]=-20;
sine[5418]=-20;
sine[5419]=-20;
sine[5420]=-20;
sine[5421]=-20;
sine[5422]=-20;
sine[5423]=-21;
sine[5424]=-21;
sine[5425]=-21;
sine[5426]=-21;
sine[5427]=-21;
sine[5428]=-21;
sine[5429]=-21;
sine[5430]=-21;
sine[5431]=-21;
sine[5432]=-21;
sine[5433]=-21;
sine[5434]=-21;
sine[5435]=-21;
sine[5436]=-21;
sine[5437]=-21;
sine[5438]=-21;
sine[5439]=-21;
sine[5440]=-21;
sine[5441]=-21;
sine[5442]=-21;
sine[5443]=-21;
sine[5444]=-22;
sine[5445]=-22;
sine[5446]=-22;
sine[5447]=-22;
sine[5448]=-22;
sine[5449]=-22;
sine[5450]=-22;
sine[5451]=-22;
sine[5452]=-22;
sine[5453]=-22;
sine[5454]=-22;
sine[5455]=-22;
sine[5456]=-22;
sine[5457]=-22;
sine[5458]=-22;
sine[5459]=-22;
sine[5460]=-22;
sine[5461]=-22;
sine[5462]=-22;
sine[5463]=-22;
sine[5464]=-22;
sine[5465]=-23;
sine[5466]=-23;
sine[5467]=-23;
sine[5468]=-23;
sine[5469]=-23;
sine[5470]=-23;
sine[5471]=-23;
sine[5472]=-23;
sine[5473]=-23;
sine[5474]=-23;
sine[5475]=-23;
sine[5476]=-23;
sine[5477]=-23;
sine[5478]=-23;
sine[5479]=-23;
sine[5480]=-23;
sine[5481]=-23;
sine[5482]=-23;
sine[5483]=-23;
sine[5484]=-23;
sine[5485]=-23;
sine[5486]=-23;
sine[5487]=-24;
sine[5488]=-24;
sine[5489]=-24;
sine[5490]=-24;
sine[5491]=-24;
sine[5492]=-24;
sine[5493]=-24;
sine[5494]=-24;
sine[5495]=-24;
sine[5496]=-24;
sine[5497]=-24;
sine[5498]=-24;
sine[5499]=-24;
sine[5500]=-24;
sine[5501]=-24;
sine[5502]=-24;
sine[5503]=-24;
sine[5504]=-24;
sine[5505]=-24;
sine[5506]=-24;
sine[5507]=-24;
sine[5508]=-25;
sine[5509]=-25;
sine[5510]=-25;
sine[5511]=-25;
sine[5512]=-25;
sine[5513]=-25;
sine[5514]=-25;
sine[5515]=-25;
sine[5516]=-25;
sine[5517]=-25;
sine[5518]=-25;
sine[5519]=-25;
sine[5520]=-25;
sine[5521]=-25;
sine[5522]=-25;
sine[5523]=-25;
sine[5524]=-25;
sine[5525]=-25;
sine[5526]=-25;
sine[5527]=-25;
sine[5528]=-25;
sine[5529]=-25;
sine[5530]=-26;
sine[5531]=-26;
sine[5532]=-26;
sine[5533]=-26;
sine[5534]=-26;
sine[5535]=-26;
sine[5536]=-26;
sine[5537]=-26;
sine[5538]=-26;
sine[5539]=-26;
sine[5540]=-26;
sine[5541]=-26;
sine[5542]=-26;
sine[5543]=-26;
sine[5544]=-26;
sine[5545]=-26;
sine[5546]=-26;
sine[5547]=-26;
sine[5548]=-26;
sine[5549]=-26;
sine[5550]=-26;
sine[5551]=-27;
sine[5552]=-27;
sine[5553]=-27;
sine[5554]=-27;
sine[5555]=-27;
sine[5556]=-27;
sine[5557]=-27;
sine[5558]=-27;
sine[5559]=-27;
sine[5560]=-27;
sine[5561]=-27;
sine[5562]=-27;
sine[5563]=-27;
sine[5564]=-27;
sine[5565]=-27;
sine[5566]=-27;
sine[5567]=-27;
sine[5568]=-27;
sine[5569]=-27;
sine[5570]=-27;
sine[5571]=-27;
sine[5572]=-27;
sine[5573]=-28;
sine[5574]=-28;
sine[5575]=-28;
sine[5576]=-28;
sine[5577]=-28;
sine[5578]=-28;
sine[5579]=-28;
sine[5580]=-28;
sine[5581]=-28;
sine[5582]=-28;
sine[5583]=-28;
sine[5584]=-28;
sine[5585]=-28;
sine[5586]=-28;
sine[5587]=-28;
sine[5588]=-28;
sine[5589]=-28;
sine[5590]=-28;
sine[5591]=-28;
sine[5592]=-28;
sine[5593]=-28;
sine[5594]=-28;
sine[5595]=-29;
sine[5596]=-29;
sine[5597]=-29;
sine[5598]=-29;
sine[5599]=-29;
sine[5600]=-29;
sine[5601]=-29;
sine[5602]=-29;
sine[5603]=-29;
sine[5604]=-29;
sine[5605]=-29;
sine[5606]=-29;
sine[5607]=-29;
sine[5608]=-29;
sine[5609]=-29;
sine[5610]=-29;
sine[5611]=-29;
sine[5612]=-29;
sine[5613]=-29;
sine[5614]=-29;
sine[5615]=-29;
sine[5616]=-29;
sine[5617]=-30;
sine[5618]=-30;
sine[5619]=-30;
sine[5620]=-30;
sine[5621]=-30;
sine[5622]=-30;
sine[5623]=-30;
sine[5624]=-30;
sine[5625]=-30;
sine[5626]=-30;
sine[5627]=-30;
sine[5628]=-30;
sine[5629]=-30;
sine[5630]=-30;
sine[5631]=-30;
sine[5632]=-30;
sine[5633]=-30;
sine[5634]=-30;
sine[5635]=-30;
sine[5636]=-30;
sine[5637]=-30;
sine[5638]=-30;
sine[5639]=-31;
sine[5640]=-31;
sine[5641]=-31;
sine[5642]=-31;
sine[5643]=-31;
sine[5644]=-31;
sine[5645]=-31;
sine[5646]=-31;
sine[5647]=-31;
sine[5648]=-31;
sine[5649]=-31;
sine[5650]=-31;
sine[5651]=-31;
sine[5652]=-31;
sine[5653]=-31;
sine[5654]=-31;
sine[5655]=-31;
sine[5656]=-31;
sine[5657]=-31;
sine[5658]=-31;
sine[5659]=-31;
sine[5660]=-31;
sine[5661]=-32;
sine[5662]=-32;
sine[5663]=-32;
sine[5664]=-32;
sine[5665]=-32;
sine[5666]=-32;
sine[5667]=-32;
sine[5668]=-32;
sine[5669]=-32;
sine[5670]=-32;
sine[5671]=-32;
sine[5672]=-32;
sine[5673]=-32;
sine[5674]=-32;
sine[5675]=-32;
sine[5676]=-32;
sine[5677]=-32;
sine[5678]=-32;
sine[5679]=-32;
sine[5680]=-32;
sine[5681]=-32;
sine[5682]=-32;
sine[5683]=-33;
sine[5684]=-33;
sine[5685]=-33;
sine[5686]=-33;
sine[5687]=-33;
sine[5688]=-33;
sine[5689]=-33;
sine[5690]=-33;
sine[5691]=-33;
sine[5692]=-33;
sine[5693]=-33;
sine[5694]=-33;
sine[5695]=-33;
sine[5696]=-33;
sine[5697]=-33;
sine[5698]=-33;
sine[5699]=-33;
sine[5700]=-33;
sine[5701]=-33;
sine[5702]=-33;
sine[5703]=-33;
sine[5704]=-33;
sine[5705]=-33;
sine[5706]=-34;
sine[5707]=-34;
sine[5708]=-34;
sine[5709]=-34;
sine[5710]=-34;
sine[5711]=-34;
sine[5712]=-34;
sine[5713]=-34;
sine[5714]=-34;
sine[5715]=-34;
sine[5716]=-34;
sine[5717]=-34;
sine[5718]=-34;
sine[5719]=-34;
sine[5720]=-34;
sine[5721]=-34;
sine[5722]=-34;
sine[5723]=-34;
sine[5724]=-34;
sine[5725]=-34;
sine[5726]=-34;
sine[5727]=-34;
sine[5728]=-35;
sine[5729]=-35;
sine[5730]=-35;
sine[5731]=-35;
sine[5732]=-35;
sine[5733]=-35;
sine[5734]=-35;
sine[5735]=-35;
sine[5736]=-35;
sine[5737]=-35;
sine[5738]=-35;
sine[5739]=-35;
sine[5740]=-35;
sine[5741]=-35;
sine[5742]=-35;
sine[5743]=-35;
sine[5744]=-35;
sine[5745]=-35;
sine[5746]=-35;
sine[5747]=-35;
sine[5748]=-35;
sine[5749]=-35;
sine[5750]=-35;
sine[5751]=-36;
sine[5752]=-36;
sine[5753]=-36;
sine[5754]=-36;
sine[5755]=-36;
sine[5756]=-36;
sine[5757]=-36;
sine[5758]=-36;
sine[5759]=-36;
sine[5760]=-36;
sine[5761]=-36;
sine[5762]=-36;
sine[5763]=-36;
sine[5764]=-36;
sine[5765]=-36;
sine[5766]=-36;
sine[5767]=-36;
sine[5768]=-36;
sine[5769]=-36;
sine[5770]=-36;
sine[5771]=-36;
sine[5772]=-36;
sine[5773]=-36;
sine[5774]=-37;
sine[5775]=-37;
sine[5776]=-37;
sine[5777]=-37;
sine[5778]=-37;
sine[5779]=-37;
sine[5780]=-37;
sine[5781]=-37;
sine[5782]=-37;
sine[5783]=-37;
sine[5784]=-37;
sine[5785]=-37;
sine[5786]=-37;
sine[5787]=-37;
sine[5788]=-37;
sine[5789]=-37;
sine[5790]=-37;
sine[5791]=-37;
sine[5792]=-37;
sine[5793]=-37;
sine[5794]=-37;
sine[5795]=-37;
sine[5796]=-37;
sine[5797]=-38;
sine[5798]=-38;
sine[5799]=-38;
sine[5800]=-38;
sine[5801]=-38;
sine[5802]=-38;
sine[5803]=-38;
sine[5804]=-38;
sine[5805]=-38;
sine[5806]=-38;
sine[5807]=-38;
sine[5808]=-38;
sine[5809]=-38;
sine[5810]=-38;
sine[5811]=-38;
sine[5812]=-38;
sine[5813]=-38;
sine[5814]=-38;
sine[5815]=-38;
sine[5816]=-38;
sine[5817]=-38;
sine[5818]=-38;
sine[5819]=-38;
sine[5820]=-38;
sine[5821]=-39;
sine[5822]=-39;
sine[5823]=-39;
sine[5824]=-39;
sine[5825]=-39;
sine[5826]=-39;
sine[5827]=-39;
sine[5828]=-39;
sine[5829]=-39;
sine[5830]=-39;
sine[5831]=-39;
sine[5832]=-39;
sine[5833]=-39;
sine[5834]=-39;
sine[5835]=-39;
sine[5836]=-39;
sine[5837]=-39;
sine[5838]=-39;
sine[5839]=-39;
sine[5840]=-39;
sine[5841]=-39;
sine[5842]=-39;
sine[5843]=-39;
sine[5844]=-40;
sine[5845]=-40;
sine[5846]=-40;
sine[5847]=-40;
sine[5848]=-40;
sine[5849]=-40;
sine[5850]=-40;
sine[5851]=-40;
sine[5852]=-40;
sine[5853]=-40;
sine[5854]=-40;
sine[5855]=-40;
sine[5856]=-40;
sine[5857]=-40;
sine[5858]=-40;
sine[5859]=-40;
sine[5860]=-40;
sine[5861]=-40;
sine[5862]=-40;
sine[5863]=-40;
sine[5864]=-40;
sine[5865]=-40;
sine[5866]=-40;
sine[5867]=-40;
sine[5868]=-41;
sine[5869]=-41;
sine[5870]=-41;
sine[5871]=-41;
sine[5872]=-41;
sine[5873]=-41;
sine[5874]=-41;
sine[5875]=-41;
sine[5876]=-41;
sine[5877]=-41;
sine[5878]=-41;
sine[5879]=-41;
sine[5880]=-41;
sine[5881]=-41;
sine[5882]=-41;
sine[5883]=-41;
sine[5884]=-41;
sine[5885]=-41;
sine[5886]=-41;
sine[5887]=-41;
sine[5888]=-41;
sine[5889]=-41;
sine[5890]=-41;
sine[5891]=-41;
sine[5892]=-42;
sine[5893]=-42;
sine[5894]=-42;
sine[5895]=-42;
sine[5896]=-42;
sine[5897]=-42;
sine[5898]=-42;
sine[5899]=-42;
sine[5900]=-42;
sine[5901]=-42;
sine[5902]=-42;
sine[5903]=-42;
sine[5904]=-42;
sine[5905]=-42;
sine[5906]=-42;
sine[5907]=-42;
sine[5908]=-42;
sine[5909]=-42;
sine[5910]=-42;
sine[5911]=-42;
sine[5912]=-42;
sine[5913]=-42;
sine[5914]=-42;
sine[5915]=-42;
sine[5916]=-43;
sine[5917]=-43;
sine[5918]=-43;
sine[5919]=-43;
sine[5920]=-43;
sine[5921]=-43;
sine[5922]=-43;
sine[5923]=-43;
sine[5924]=-43;
sine[5925]=-43;
sine[5926]=-43;
sine[5927]=-43;
sine[5928]=-43;
sine[5929]=-43;
sine[5930]=-43;
sine[5931]=-43;
sine[5932]=-43;
sine[5933]=-43;
sine[5934]=-43;
sine[5935]=-43;
sine[5936]=-43;
sine[5937]=-43;
sine[5938]=-43;
sine[5939]=-43;
sine[5940]=-44;
sine[5941]=-44;
sine[5942]=-44;
sine[5943]=-44;
sine[5944]=-44;
sine[5945]=-44;
sine[5946]=-44;
sine[5947]=-44;
sine[5948]=-44;
sine[5949]=-44;
sine[5950]=-44;
sine[5951]=-44;
sine[5952]=-44;
sine[5953]=-44;
sine[5954]=-44;
sine[5955]=-44;
sine[5956]=-44;
sine[5957]=-44;
sine[5958]=-44;
sine[5959]=-44;
sine[5960]=-44;
sine[5961]=-44;
sine[5962]=-44;
sine[5963]=-44;
sine[5964]=-44;
sine[5965]=-45;
sine[5966]=-45;
sine[5967]=-45;
sine[5968]=-45;
sine[5969]=-45;
sine[5970]=-45;
sine[5971]=-45;
sine[5972]=-45;
sine[5973]=-45;
sine[5974]=-45;
sine[5975]=-45;
sine[5976]=-45;
sine[5977]=-45;
sine[5978]=-45;
sine[5979]=-45;
sine[5980]=-45;
sine[5981]=-45;
sine[5982]=-45;
sine[5983]=-45;
sine[5984]=-45;
sine[5985]=-45;
sine[5986]=-45;
sine[5987]=-45;
sine[5988]=-45;
sine[5989]=-45;
sine[5990]=-46;
sine[5991]=-46;
sine[5992]=-46;
sine[5993]=-46;
sine[5994]=-46;
sine[5995]=-46;
sine[5996]=-46;
sine[5997]=-46;
sine[5998]=-46;
sine[5999]=-46;
sine[6000]=-46;
sine[6001]=-46;
sine[6002]=-46;
sine[6003]=-46;
sine[6004]=-46;
sine[6005]=-46;
sine[6006]=-46;
sine[6007]=-46;
sine[6008]=-46;
sine[6009]=-46;
sine[6010]=-46;
sine[6011]=-46;
sine[6012]=-46;
sine[6013]=-46;
sine[6014]=-46;
sine[6015]=-47;
sine[6016]=-47;
sine[6017]=-47;
sine[6018]=-47;
sine[6019]=-47;
sine[6020]=-47;
sine[6021]=-47;
sine[6022]=-47;
sine[6023]=-47;
sine[6024]=-47;
sine[6025]=-47;
sine[6026]=-47;
sine[6027]=-47;
sine[6028]=-47;
sine[6029]=-47;
sine[6030]=-47;
sine[6031]=-47;
sine[6032]=-47;
sine[6033]=-47;
sine[6034]=-47;
sine[6035]=-47;
sine[6036]=-47;
sine[6037]=-47;
sine[6038]=-47;
sine[6039]=-47;
sine[6040]=-47;
sine[6041]=-48;
sine[6042]=-48;
sine[6043]=-48;
sine[6044]=-48;
sine[6045]=-48;
sine[6046]=-48;
sine[6047]=-48;
sine[6048]=-48;
sine[6049]=-48;
sine[6050]=-48;
sine[6051]=-48;
sine[6052]=-48;
sine[6053]=-48;
sine[6054]=-48;
sine[6055]=-48;
sine[6056]=-48;
sine[6057]=-48;
sine[6058]=-48;
sine[6059]=-48;
sine[6060]=-48;
sine[6061]=-48;
sine[6062]=-48;
sine[6063]=-48;
sine[6064]=-48;
sine[6065]=-48;
sine[6066]=-49;
sine[6067]=-49;
sine[6068]=-49;
sine[6069]=-49;
sine[6070]=-49;
sine[6071]=-49;
sine[6072]=-49;
sine[6073]=-49;
sine[6074]=-49;
sine[6075]=-49;
sine[6076]=-49;
sine[6077]=-49;
sine[6078]=-49;
sine[6079]=-49;
sine[6080]=-49;
sine[6081]=-49;
sine[6082]=-49;
sine[6083]=-49;
sine[6084]=-49;
sine[6085]=-49;
sine[6086]=-49;
sine[6087]=-49;
sine[6088]=-49;
sine[6089]=-49;
sine[6090]=-49;
sine[6091]=-49;
sine[6092]=-49;
sine[6093]=-50;
sine[6094]=-50;
sine[6095]=-50;
sine[6096]=-50;
sine[6097]=-50;
sine[6098]=-50;
sine[6099]=-50;
sine[6100]=-50;
sine[6101]=-50;
sine[6102]=-50;
sine[6103]=-50;
sine[6104]=-50;
sine[6105]=-50;
sine[6106]=-50;
sine[6107]=-50;
sine[6108]=-50;
sine[6109]=-50;
sine[6110]=-50;
sine[6111]=-50;
sine[6112]=-50;
sine[6113]=-50;
sine[6114]=-50;
sine[6115]=-50;
sine[6116]=-50;
sine[6117]=-50;
sine[6118]=-50;
sine[6119]=-51;
sine[6120]=-51;
sine[6121]=-51;
sine[6122]=-51;
sine[6123]=-51;
sine[6124]=-51;
sine[6125]=-51;
sine[6126]=-51;
sine[6127]=-51;
sine[6128]=-51;
sine[6129]=-51;
sine[6130]=-51;
sine[6131]=-51;
sine[6132]=-51;
sine[6133]=-51;
sine[6134]=-51;
sine[6135]=-51;
sine[6136]=-51;
sine[6137]=-51;
sine[6138]=-51;
sine[6139]=-51;
sine[6140]=-51;
sine[6141]=-51;
sine[6142]=-51;
sine[6143]=-51;
sine[6144]=-51;
sine[6145]=-51;
sine[6146]=-52;
sine[6147]=-52;
sine[6148]=-52;
sine[6149]=-52;
sine[6150]=-52;
sine[6151]=-52;
sine[6152]=-52;
sine[6153]=-52;
sine[6154]=-52;
sine[6155]=-52;
sine[6156]=-52;
sine[6157]=-52;
sine[6158]=-52;
sine[6159]=-52;
sine[6160]=-52;
sine[6161]=-52;
sine[6162]=-52;
sine[6163]=-52;
sine[6164]=-52;
sine[6165]=-52;
sine[6166]=-52;
sine[6167]=-52;
sine[6168]=-52;
sine[6169]=-52;
sine[6170]=-52;
sine[6171]=-52;
sine[6172]=-52;
sine[6173]=-53;
sine[6174]=-53;
sine[6175]=-53;
sine[6176]=-53;
sine[6177]=-53;
sine[6178]=-53;
sine[6179]=-53;
sine[6180]=-53;
sine[6181]=-53;
sine[6182]=-53;
sine[6183]=-53;
sine[6184]=-53;
sine[6185]=-53;
sine[6186]=-53;
sine[6187]=-53;
sine[6188]=-53;
sine[6189]=-53;
sine[6190]=-53;
sine[6191]=-53;
sine[6192]=-53;
sine[6193]=-53;
sine[6194]=-53;
sine[6195]=-53;
sine[6196]=-53;
sine[6197]=-53;
sine[6198]=-53;
sine[6199]=-53;
sine[6200]=-53;
sine[6201]=-54;
sine[6202]=-54;
sine[6203]=-54;
sine[6204]=-54;
sine[6205]=-54;
sine[6206]=-54;
sine[6207]=-54;
sine[6208]=-54;
sine[6209]=-54;
sine[6210]=-54;
sine[6211]=-54;
sine[6212]=-54;
sine[6213]=-54;
sine[6214]=-54;
sine[6215]=-54;
sine[6216]=-54;
sine[6217]=-54;
sine[6218]=-54;
sine[6219]=-54;
sine[6220]=-54;
sine[6221]=-54;
sine[6222]=-54;
sine[6223]=-54;
sine[6224]=-54;
sine[6225]=-54;
sine[6226]=-54;
sine[6227]=-54;
sine[6228]=-54;
sine[6229]=-55;
sine[6230]=-55;
sine[6231]=-55;
sine[6232]=-55;
sine[6233]=-55;
sine[6234]=-55;
sine[6235]=-55;
sine[6236]=-55;
sine[6237]=-55;
sine[6238]=-55;
sine[6239]=-55;
sine[6240]=-55;
sine[6241]=-55;
sine[6242]=-55;
sine[6243]=-55;
sine[6244]=-55;
sine[6245]=-55;
sine[6246]=-55;
sine[6247]=-55;
sine[6248]=-55;
sine[6249]=-55;
sine[6250]=-55;
sine[6251]=-55;
sine[6252]=-55;
sine[6253]=-55;
sine[6254]=-55;
sine[6255]=-55;
sine[6256]=-55;
sine[6257]=-55;
sine[6258]=-56;
sine[6259]=-56;
sine[6260]=-56;
sine[6261]=-56;
sine[6262]=-56;
sine[6263]=-56;
sine[6264]=-56;
sine[6265]=-56;
sine[6266]=-56;
sine[6267]=-56;
sine[6268]=-56;
sine[6269]=-56;
sine[6270]=-56;
sine[6271]=-56;
sine[6272]=-56;
sine[6273]=-56;
sine[6274]=-56;
sine[6275]=-56;
sine[6276]=-56;
sine[6277]=-56;
sine[6278]=-56;
sine[6279]=-56;
sine[6280]=-56;
sine[6281]=-56;
sine[6282]=-56;
sine[6283]=-56;
sine[6284]=-56;
sine[6285]=-56;
sine[6286]=-56;
sine[6287]=-57;
sine[6288]=-57;
sine[6289]=-57;
sine[6290]=-57;
sine[6291]=-57;
sine[6292]=-57;
sine[6293]=-57;
sine[6294]=-57;
sine[6295]=-57;
sine[6296]=-57;
sine[6297]=-57;
sine[6298]=-57;
sine[6299]=-57;
sine[6300]=-57;
sine[6301]=-57;
sine[6302]=-57;
sine[6303]=-57;
sine[6304]=-57;
sine[6305]=-57;
sine[6306]=-57;
sine[6307]=-57;
sine[6308]=-57;
sine[6309]=-57;
sine[6310]=-57;
sine[6311]=-57;
sine[6312]=-57;
sine[6313]=-57;
sine[6314]=-57;
sine[6315]=-57;
sine[6316]=-57;
sine[6317]=-58;
sine[6318]=-58;
sine[6319]=-58;
sine[6320]=-58;
sine[6321]=-58;
sine[6322]=-58;
sine[6323]=-58;
sine[6324]=-58;
sine[6325]=-58;
sine[6326]=-58;
sine[6327]=-58;
sine[6328]=-58;
sine[6329]=-58;
sine[6330]=-58;
sine[6331]=-58;
sine[6332]=-58;
sine[6333]=-58;
sine[6334]=-58;
sine[6335]=-58;
sine[6336]=-58;
sine[6337]=-58;
sine[6338]=-58;
sine[6339]=-58;
sine[6340]=-58;
sine[6341]=-58;
sine[6342]=-58;
sine[6343]=-58;
sine[6344]=-58;
sine[6345]=-58;
sine[6346]=-58;
sine[6347]=-59;
sine[6348]=-59;
sine[6349]=-59;
sine[6350]=-59;
sine[6351]=-59;
sine[6352]=-59;
sine[6353]=-59;
sine[6354]=-59;
sine[6355]=-59;
sine[6356]=-59;
sine[6357]=-59;
sine[6358]=-59;
sine[6359]=-59;
sine[6360]=-59;
sine[6361]=-59;
sine[6362]=-59;
sine[6363]=-59;
sine[6364]=-59;
sine[6365]=-59;
sine[6366]=-59;
sine[6367]=-59;
sine[6368]=-59;
sine[6369]=-59;
sine[6370]=-59;
sine[6371]=-59;
sine[6372]=-59;
sine[6373]=-59;
sine[6374]=-59;
sine[6375]=-59;
sine[6376]=-59;
sine[6377]=-59;
sine[6378]=-60;
sine[6379]=-60;
sine[6380]=-60;
sine[6381]=-60;
sine[6382]=-60;
sine[6383]=-60;
sine[6384]=-60;
sine[6385]=-60;
sine[6386]=-60;
sine[6387]=-60;
sine[6388]=-60;
sine[6389]=-60;
sine[6390]=-60;
sine[6391]=-60;
sine[6392]=-60;
sine[6393]=-60;
sine[6394]=-60;
sine[6395]=-60;
sine[6396]=-60;
sine[6397]=-60;
sine[6398]=-60;
sine[6399]=-60;
sine[6400]=-60;
sine[6401]=-60;
sine[6402]=-60;
sine[6403]=-60;
sine[6404]=-60;
sine[6405]=-60;
sine[6406]=-60;
sine[6407]=-60;
sine[6408]=-60;
sine[6409]=-60;
sine[6410]=-61;
sine[6411]=-61;
sine[6412]=-61;
sine[6413]=-61;
sine[6414]=-61;
sine[6415]=-61;
sine[6416]=-61;
sine[6417]=-61;
sine[6418]=-61;
sine[6419]=-61;
sine[6420]=-61;
sine[6421]=-61;
sine[6422]=-61;
sine[6423]=-61;
sine[6424]=-61;
sine[6425]=-61;
sine[6426]=-61;
sine[6427]=-61;
sine[6428]=-61;
sine[6429]=-61;
sine[6430]=-61;
sine[6431]=-61;
sine[6432]=-61;
sine[6433]=-61;
sine[6434]=-61;
sine[6435]=-61;
sine[6436]=-61;
sine[6437]=-61;
sine[6438]=-61;
sine[6439]=-61;
sine[6440]=-61;
sine[6441]=-61;
sine[6442]=-61;
sine[6443]=-62;
sine[6444]=-62;
sine[6445]=-62;
sine[6446]=-62;
sine[6447]=-62;
sine[6448]=-62;
sine[6449]=-62;
sine[6450]=-62;
sine[6451]=-62;
sine[6452]=-62;
sine[6453]=-62;
sine[6454]=-62;
sine[6455]=-62;
sine[6456]=-62;
sine[6457]=-62;
sine[6458]=-62;
sine[6459]=-62;
sine[6460]=-62;
sine[6461]=-62;
sine[6462]=-62;
sine[6463]=-62;
sine[6464]=-62;
sine[6465]=-62;
sine[6466]=-62;
sine[6467]=-62;
sine[6468]=-62;
sine[6469]=-62;
sine[6470]=-62;
sine[6471]=-62;
sine[6472]=-62;
sine[6473]=-62;
sine[6474]=-62;
sine[6475]=-62;
sine[6476]=-63;
sine[6477]=-63;
sine[6478]=-63;
sine[6479]=-63;
sine[6480]=-63;
sine[6481]=-63;
sine[6482]=-63;
sine[6483]=-63;
sine[6484]=-63;
sine[6485]=-63;
sine[6486]=-63;
sine[6487]=-63;
sine[6488]=-63;
sine[6489]=-63;
sine[6490]=-63;
sine[6491]=-63;
sine[6492]=-63;
sine[6493]=-63;
sine[6494]=-63;
sine[6495]=-63;
sine[6496]=-63;
sine[6497]=-63;
sine[6498]=-63;
sine[6499]=-63;
sine[6500]=-63;
sine[6501]=-63;
sine[6502]=-63;
sine[6503]=-63;
sine[6504]=-63;
sine[6505]=-63;
sine[6506]=-63;
sine[6507]=-63;
sine[6508]=-63;
sine[6509]=-63;
sine[6510]=-63;
sine[6511]=-64;
sine[6512]=-64;
sine[6513]=-64;
sine[6514]=-64;
sine[6515]=-64;
sine[6516]=-64;
sine[6517]=-64;
sine[6518]=-64;
sine[6519]=-64;
sine[6520]=-64;
sine[6521]=-64;
sine[6522]=-64;
sine[6523]=-64;
sine[6524]=-64;
sine[6525]=-64;
sine[6526]=-64;
sine[6527]=-64;
sine[6528]=-64;
sine[6529]=-64;
sine[6530]=-64;
sine[6531]=-64;
sine[6532]=-64;
sine[6533]=-64;
sine[6534]=-64;
sine[6535]=-64;
sine[6536]=-64;
sine[6537]=-64;
sine[6538]=-64;
sine[6539]=-64;
sine[6540]=-64;
sine[6541]=-64;
sine[6542]=-64;
sine[6543]=-64;
sine[6544]=-64;
sine[6545]=-64;
sine[6546]=-65;
sine[6547]=-65;
sine[6548]=-65;
sine[6549]=-65;
sine[6550]=-65;
sine[6551]=-65;
sine[6552]=-65;
sine[6553]=-65;
sine[6554]=-65;
sine[6555]=-65;
sine[6556]=-65;
sine[6557]=-65;
sine[6558]=-65;
sine[6559]=-65;
sine[6560]=-65;
sine[6561]=-65;
sine[6562]=-65;
sine[6563]=-65;
sine[6564]=-65;
sine[6565]=-65;
sine[6566]=-65;
sine[6567]=-65;
sine[6568]=-65;
sine[6569]=-65;
sine[6570]=-65;
sine[6571]=-65;
sine[6572]=-65;
sine[6573]=-65;
sine[6574]=-65;
sine[6575]=-65;
sine[6576]=-65;
sine[6577]=-65;
sine[6578]=-65;
sine[6579]=-65;
sine[6580]=-65;
sine[6581]=-65;
sine[6582]=-65;
sine[6583]=-66;
sine[6584]=-66;
sine[6585]=-66;
sine[6586]=-66;
sine[6587]=-66;
sine[6588]=-66;
sine[6589]=-66;
sine[6590]=-66;
sine[6591]=-66;
sine[6592]=-66;
sine[6593]=-66;
sine[6594]=-66;
sine[6595]=-66;
sine[6596]=-66;
sine[6597]=-66;
sine[6598]=-66;
sine[6599]=-66;
sine[6600]=-66;
sine[6601]=-66;
sine[6602]=-66;
sine[6603]=-66;
sine[6604]=-66;
sine[6605]=-66;
sine[6606]=-66;
sine[6607]=-66;
sine[6608]=-66;
sine[6609]=-66;
sine[6610]=-66;
sine[6611]=-66;
sine[6612]=-66;
sine[6613]=-66;
sine[6614]=-66;
sine[6615]=-66;
sine[6616]=-66;
sine[6617]=-66;
sine[6618]=-66;
sine[6619]=-66;
sine[6620]=-66;
sine[6621]=-67;
sine[6622]=-67;
sine[6623]=-67;
sine[6624]=-67;
sine[6625]=-67;
sine[6626]=-67;
sine[6627]=-67;
sine[6628]=-67;
sine[6629]=-67;
sine[6630]=-67;
sine[6631]=-67;
sine[6632]=-67;
sine[6633]=-67;
sine[6634]=-67;
sine[6635]=-67;
sine[6636]=-67;
sine[6637]=-67;
sine[6638]=-67;
sine[6639]=-67;
sine[6640]=-67;
sine[6641]=-67;
sine[6642]=-67;
sine[6643]=-67;
sine[6644]=-67;
sine[6645]=-67;
sine[6646]=-67;
sine[6647]=-67;
sine[6648]=-67;
sine[6649]=-67;
sine[6650]=-67;
sine[6651]=-67;
sine[6652]=-67;
sine[6653]=-67;
sine[6654]=-67;
sine[6655]=-67;
sine[6656]=-67;
sine[6657]=-67;
sine[6658]=-67;
sine[6659]=-67;
sine[6660]=-67;
sine[6661]=-68;
sine[6662]=-68;
sine[6663]=-68;
sine[6664]=-68;
sine[6665]=-68;
sine[6666]=-68;
sine[6667]=-68;
sine[6668]=-68;
sine[6669]=-68;
sine[6670]=-68;
sine[6671]=-68;
sine[6672]=-68;
sine[6673]=-68;
sine[6674]=-68;
sine[6675]=-68;
sine[6676]=-68;
sine[6677]=-68;
sine[6678]=-68;
sine[6679]=-68;
sine[6680]=-68;
sine[6681]=-68;
sine[6682]=-68;
sine[6683]=-68;
sine[6684]=-68;
sine[6685]=-68;
sine[6686]=-68;
sine[6687]=-68;
sine[6688]=-68;
sine[6689]=-68;
sine[6690]=-68;
sine[6691]=-68;
sine[6692]=-68;
sine[6693]=-68;
sine[6694]=-68;
sine[6695]=-68;
sine[6696]=-68;
sine[6697]=-68;
sine[6698]=-68;
sine[6699]=-68;
sine[6700]=-68;
sine[6701]=-68;
sine[6702]=-69;
sine[6703]=-69;
sine[6704]=-69;
sine[6705]=-69;
sine[6706]=-69;
sine[6707]=-69;
sine[6708]=-69;
sine[6709]=-69;
sine[6710]=-69;
sine[6711]=-69;
sine[6712]=-69;
sine[6713]=-69;
sine[6714]=-69;
sine[6715]=-69;
sine[6716]=-69;
sine[6717]=-69;
sine[6718]=-69;
sine[6719]=-69;
sine[6720]=-69;
sine[6721]=-69;
sine[6722]=-69;
sine[6723]=-69;
sine[6724]=-69;
sine[6725]=-69;
sine[6726]=-69;
sine[6727]=-69;
sine[6728]=-69;
sine[6729]=-69;
sine[6730]=-69;
sine[6731]=-69;
sine[6732]=-69;
sine[6733]=-69;
sine[6734]=-69;
sine[6735]=-69;
sine[6736]=-69;
sine[6737]=-69;
sine[6738]=-69;
sine[6739]=-69;
sine[6740]=-69;
sine[6741]=-69;
sine[6742]=-69;
sine[6743]=-69;
sine[6744]=-69;
sine[6745]=-69;
sine[6746]=-70;
sine[6747]=-70;
sine[6748]=-70;
sine[6749]=-70;
sine[6750]=-70;
sine[6751]=-70;
sine[6752]=-70;
sine[6753]=-70;
sine[6754]=-70;
sine[6755]=-70;
sine[6756]=-70;
sine[6757]=-70;
sine[6758]=-70;
sine[6759]=-70;
sine[6760]=-70;
sine[6761]=-70;
sine[6762]=-70;
sine[6763]=-70;
sine[6764]=-70;
sine[6765]=-70;
sine[6766]=-70;
sine[6767]=-70;
sine[6768]=-70;
sine[6769]=-70;
sine[6770]=-70;
sine[6771]=-70;
sine[6772]=-70;
sine[6773]=-70;
sine[6774]=-70;
sine[6775]=-70;
sine[6776]=-70;
sine[6777]=-70;
sine[6778]=-70;
sine[6779]=-70;
sine[6780]=-70;
sine[6781]=-70;
sine[6782]=-70;
sine[6783]=-70;
sine[6784]=-70;
sine[6785]=-70;
sine[6786]=-70;
sine[6787]=-70;
sine[6788]=-70;
sine[6789]=-70;
sine[6790]=-70;
sine[6791]=-71;
sine[6792]=-71;
sine[6793]=-71;
sine[6794]=-71;
sine[6795]=-71;
sine[6796]=-71;
sine[6797]=-71;
sine[6798]=-71;
sine[6799]=-71;
sine[6800]=-71;
sine[6801]=-71;
sine[6802]=-71;
sine[6803]=-71;
sine[6804]=-71;
sine[6805]=-71;
sine[6806]=-71;
sine[6807]=-71;
sine[6808]=-71;
sine[6809]=-71;
sine[6810]=-71;
sine[6811]=-71;
sine[6812]=-71;
sine[6813]=-71;
sine[6814]=-71;
sine[6815]=-71;
sine[6816]=-71;
sine[6817]=-71;
sine[6818]=-71;
sine[6819]=-71;
sine[6820]=-71;
sine[6821]=-71;
sine[6822]=-71;
sine[6823]=-71;
sine[6824]=-71;
sine[6825]=-71;
sine[6826]=-71;
sine[6827]=-71;
sine[6828]=-71;
sine[6829]=-71;
sine[6830]=-71;
sine[6831]=-71;
sine[6832]=-71;
sine[6833]=-71;
sine[6834]=-71;
sine[6835]=-71;
sine[6836]=-71;
sine[6837]=-71;
sine[6838]=-71;
sine[6839]=-71;
sine[6840]=-72;
sine[6841]=-72;
sine[6842]=-72;
sine[6843]=-72;
sine[6844]=-72;
sine[6845]=-72;
sine[6846]=-72;
sine[6847]=-72;
sine[6848]=-72;
sine[6849]=-72;
sine[6850]=-72;
sine[6851]=-72;
sine[6852]=-72;
sine[6853]=-72;
sine[6854]=-72;
sine[6855]=-72;
sine[6856]=-72;
sine[6857]=-72;
sine[6858]=-72;
sine[6859]=-72;
sine[6860]=-72;
sine[6861]=-72;
sine[6862]=-72;
sine[6863]=-72;
sine[6864]=-72;
sine[6865]=-72;
sine[6866]=-72;
sine[6867]=-72;
sine[6868]=-72;
sine[6869]=-72;
sine[6870]=-72;
sine[6871]=-72;
sine[6872]=-72;
sine[6873]=-72;
sine[6874]=-72;
sine[6875]=-72;
sine[6876]=-72;
sine[6877]=-72;
sine[6878]=-72;
sine[6879]=-72;
sine[6880]=-72;
sine[6881]=-72;
sine[6882]=-72;
sine[6883]=-72;
sine[6884]=-72;
sine[6885]=-72;
sine[6886]=-72;
sine[6887]=-72;
sine[6888]=-72;
sine[6889]=-72;
sine[6890]=-72;
sine[6891]=-72;
sine[6892]=-72;
sine[6893]=-73;
sine[6894]=-73;
sine[6895]=-73;
sine[6896]=-73;
sine[6897]=-73;
sine[6898]=-73;
sine[6899]=-73;
sine[6900]=-73;
sine[6901]=-73;
sine[6902]=-73;
sine[6903]=-73;
sine[6904]=-73;
sine[6905]=-73;
sine[6906]=-73;
sine[6907]=-73;
sine[6908]=-73;
sine[6909]=-73;
sine[6910]=-73;
sine[6911]=-73;
sine[6912]=-73;
sine[6913]=-73;
sine[6914]=-73;
sine[6915]=-73;
sine[6916]=-73;
sine[6917]=-73;
sine[6918]=-73;
sine[6919]=-73;
sine[6920]=-73;
sine[6921]=-73;
sine[6922]=-73;
sine[6923]=-73;
sine[6924]=-73;
sine[6925]=-73;
sine[6926]=-73;
sine[6927]=-73;
sine[6928]=-73;
sine[6929]=-73;
sine[6930]=-73;
sine[6931]=-73;
sine[6932]=-73;
sine[6933]=-73;
sine[6934]=-73;
sine[6935]=-73;
sine[6936]=-73;
sine[6937]=-73;
sine[6938]=-73;
sine[6939]=-73;
sine[6940]=-73;
sine[6941]=-73;
sine[6942]=-73;
sine[6943]=-73;
sine[6944]=-73;
sine[6945]=-73;
sine[6946]=-73;
sine[6947]=-73;
sine[6948]=-73;
sine[6949]=-73;
sine[6950]=-74;
sine[6951]=-74;
sine[6952]=-74;
sine[6953]=-74;
sine[6954]=-74;
sine[6955]=-74;
sine[6956]=-74;
sine[6957]=-74;
sine[6958]=-74;
sine[6959]=-74;
sine[6960]=-74;
sine[6961]=-74;
sine[6962]=-74;
sine[6963]=-74;
sine[6964]=-74;
sine[6965]=-74;
sine[6966]=-74;
sine[6967]=-74;
sine[6968]=-74;
sine[6969]=-74;
sine[6970]=-74;
sine[6971]=-74;
sine[6972]=-74;
sine[6973]=-74;
sine[6974]=-74;
sine[6975]=-74;
sine[6976]=-74;
sine[6977]=-74;
sine[6978]=-74;
sine[6979]=-74;
sine[6980]=-74;
sine[6981]=-74;
sine[6982]=-74;
sine[6983]=-74;
sine[6984]=-74;
sine[6985]=-74;
sine[6986]=-74;
sine[6987]=-74;
sine[6988]=-74;
sine[6989]=-74;
sine[6990]=-74;
sine[6991]=-74;
sine[6992]=-74;
sine[6993]=-74;
sine[6994]=-74;
sine[6995]=-74;
sine[6996]=-74;
sine[6997]=-74;
sine[6998]=-74;
sine[6999]=-74;
sine[7000]=-74;
sine[7001]=-74;
sine[7002]=-74;
sine[7003]=-74;
sine[7004]=-74;
sine[7005]=-74;
sine[7006]=-74;
sine[7007]=-74;
sine[7008]=-74;
sine[7009]=-74;
sine[7010]=-74;
sine[7011]=-74;
sine[7012]=-74;
sine[7013]=-74;
sine[7014]=-75;
sine[7015]=-75;
sine[7016]=-75;
sine[7017]=-75;
sine[7018]=-75;
sine[7019]=-75;
sine[7020]=-75;
sine[7021]=-75;
sine[7022]=-75;
sine[7023]=-75;
sine[7024]=-75;
sine[7025]=-75;
sine[7026]=-75;
sine[7027]=-75;
sine[7028]=-75;
sine[7029]=-75;
sine[7030]=-75;
sine[7031]=-75;
sine[7032]=-75;
sine[7033]=-75;
sine[7034]=-75;
sine[7035]=-75;
sine[7036]=-75;
sine[7037]=-75;
sine[7038]=-75;
sine[7039]=-75;
sine[7040]=-75;
sine[7041]=-75;
sine[7042]=-75;
sine[7043]=-75;
sine[7044]=-75;
sine[7045]=-75;
sine[7046]=-75;
sine[7047]=-75;
sine[7048]=-75;
sine[7049]=-75;
sine[7050]=-75;
sine[7051]=-75;
sine[7052]=-75;
sine[7053]=-75;
sine[7054]=-75;
sine[7055]=-75;
sine[7056]=-75;
sine[7057]=-75;
sine[7058]=-75;
sine[7059]=-75;
sine[7060]=-75;
sine[7061]=-75;
sine[7062]=-75;
sine[7063]=-75;
sine[7064]=-75;
sine[7065]=-75;
sine[7066]=-75;
sine[7067]=-75;
sine[7068]=-75;
sine[7069]=-75;
sine[7070]=-75;
sine[7071]=-75;
sine[7072]=-75;
sine[7073]=-75;
sine[7074]=-75;
sine[7075]=-75;
sine[7076]=-75;
sine[7077]=-75;
sine[7078]=-75;
sine[7079]=-75;
sine[7080]=-75;
sine[7081]=-75;
sine[7082]=-75;
sine[7083]=-75;
sine[7084]=-75;
sine[7085]=-75;
sine[7086]=-75;
sine[7087]=-76;
sine[7088]=-76;
sine[7089]=-76;
sine[7090]=-76;
sine[7091]=-76;
sine[7092]=-76;
sine[7093]=-76;
sine[7094]=-76;
sine[7095]=-76;
sine[7096]=-76;
sine[7097]=-76;
sine[7098]=-76;
sine[7099]=-76;
sine[7100]=-76;
sine[7101]=-76;
sine[7102]=-76;
sine[7103]=-76;
sine[7104]=-76;
sine[7105]=-76;
sine[7106]=-76;
sine[7107]=-76;
sine[7108]=-76;
sine[7109]=-76;
sine[7110]=-76;
sine[7111]=-76;
sine[7112]=-76;
sine[7113]=-76;
sine[7114]=-76;
sine[7115]=-76;
sine[7116]=-76;
sine[7117]=-76;
sine[7118]=-76;
sine[7119]=-76;
sine[7120]=-76;
sine[7121]=-76;
sine[7122]=-76;
sine[7123]=-76;
sine[7124]=-76;
sine[7125]=-76;
sine[7126]=-76;
sine[7127]=-76;
sine[7128]=-76;
sine[7129]=-76;
sine[7130]=-76;
sine[7131]=-76;
sine[7132]=-76;
sine[7133]=-76;
sine[7134]=-76;
sine[7135]=-76;
sine[7136]=-76;
sine[7137]=-76;
sine[7138]=-76;
sine[7139]=-76;
sine[7140]=-76;
sine[7141]=-76;
sine[7142]=-76;
sine[7143]=-76;
sine[7144]=-76;
sine[7145]=-76;
sine[7146]=-76;
sine[7147]=-76;
sine[7148]=-76;
sine[7149]=-76;
sine[7150]=-76;
sine[7151]=-76;
sine[7152]=-76;
sine[7153]=-76;
sine[7154]=-76;
sine[7155]=-76;
sine[7156]=-76;
sine[7157]=-76;
sine[7158]=-76;
sine[7159]=-76;
sine[7160]=-76;
sine[7161]=-76;
sine[7162]=-76;
sine[7163]=-76;
sine[7164]=-76;
sine[7165]=-76;
sine[7166]=-76;
sine[7167]=-76;
sine[7168]=-76;
sine[7169]=-76;
sine[7170]=-76;
sine[7171]=-76;
sine[7172]=-76;
sine[7173]=-76;
sine[7174]=-76;
sine[7175]=-77;
sine[7176]=-77;
sine[7177]=-77;
sine[7178]=-77;
sine[7179]=-77;
sine[7180]=-77;
sine[7181]=-77;
sine[7182]=-77;
sine[7183]=-77;
sine[7184]=-77;
sine[7185]=-77;
sine[7186]=-77;
sine[7187]=-77;
sine[7188]=-77;
sine[7189]=-77;
sine[7190]=-77;
sine[7191]=-77;
sine[7192]=-77;
sine[7193]=-77;
sine[7194]=-77;
sine[7195]=-77;
sine[7196]=-77;
sine[7197]=-77;
sine[7198]=-77;
sine[7199]=-77;
sine[7200]=-77;
sine[7201]=-77;
sine[7202]=-77;
sine[7203]=-77;
sine[7204]=-77;
sine[7205]=-77;
sine[7206]=-77;
sine[7207]=-77;
sine[7208]=-77;
sine[7209]=-77;
sine[7210]=-77;
sine[7211]=-77;
sine[7212]=-77;
sine[7213]=-77;
sine[7214]=-77;
sine[7215]=-77;
sine[7216]=-77;
sine[7217]=-77;
sine[7218]=-77;
sine[7219]=-77;
sine[7220]=-77;
sine[7221]=-77;
sine[7222]=-77;
sine[7223]=-77;
sine[7224]=-77;
sine[7225]=-77;
sine[7226]=-77;
sine[7227]=-77;
sine[7228]=-77;
sine[7229]=-77;
sine[7230]=-77;
sine[7231]=-77;
sine[7232]=-77;
sine[7233]=-77;
sine[7234]=-77;
sine[7235]=-77;
sine[7236]=-77;
sine[7237]=-77;
sine[7238]=-77;
sine[7239]=-77;
sine[7240]=-77;
sine[7241]=-77;
sine[7242]=-77;
sine[7243]=-77;
sine[7244]=-77;
sine[7245]=-77;
sine[7246]=-77;
sine[7247]=-77;
sine[7248]=-77;
sine[7249]=-77;
sine[7250]=-77;
sine[7251]=-77;
sine[7252]=-77;
sine[7253]=-77;
sine[7254]=-77;
sine[7255]=-77;
sine[7256]=-77;
sine[7257]=-77;
sine[7258]=-77;
sine[7259]=-77;
sine[7260]=-77;
sine[7261]=-77;
sine[7262]=-77;
sine[7263]=-77;
sine[7264]=-77;
sine[7265]=-77;
sine[7266]=-77;
sine[7267]=-77;
sine[7268]=-77;
sine[7269]=-77;
sine[7270]=-77;
sine[7271]=-77;
sine[7272]=-77;
sine[7273]=-77;
sine[7274]=-77;
sine[7275]=-77;
sine[7276]=-77;
sine[7277]=-77;
sine[7278]=-77;
sine[7279]=-77;
sine[7280]=-77;
sine[7281]=-77;
sine[7282]=-77;
sine[7283]=-77;
sine[7284]=-77;
sine[7285]=-77;
sine[7286]=-77;
sine[7287]=-77;
sine[7288]=-77;
sine[7289]=-77;
sine[7290]=-77;
sine[7291]=-77;
sine[7292]=-77;
sine[7293]=-77;
sine[7294]=-77;
sine[7295]=-77;
sine[7296]=-77;
sine[7297]=-77;
sine[7298]=-77;
sine[7299]=-78;
sine[7300]=-78;
sine[7301]=-78;
sine[7302]=-78;
sine[7303]=-78;
sine[7304]=-78;
sine[7305]=-78;
sine[7306]=-78;
sine[7307]=-78;
sine[7308]=-78;
sine[7309]=-78;
sine[7310]=-78;
sine[7311]=-78;
sine[7312]=-78;
sine[7313]=-78;
sine[7314]=-78;
sine[7315]=-78;
sine[7316]=-78;
sine[7317]=-78;
sine[7318]=-78;
sine[7319]=-78;
sine[7320]=-78;
sine[7321]=-78;
sine[7322]=-78;
sine[7323]=-78;
sine[7324]=-78;
sine[7325]=-78;
sine[7326]=-78;
sine[7327]=-78;
sine[7328]=-78;
sine[7329]=-78;
sine[7330]=-78;
sine[7331]=-78;
sine[7332]=-78;
sine[7333]=-78;
sine[7334]=-78;
sine[7335]=-78;
sine[7336]=-78;
sine[7337]=-78;
sine[7338]=-78;
sine[7339]=-78;
sine[7340]=-78;
sine[7341]=-78;
sine[7342]=-78;
sine[7343]=-78;
sine[7344]=-78;
sine[7345]=-78;
sine[7346]=-78;
sine[7347]=-78;
sine[7348]=-78;
sine[7349]=-78;
sine[7350]=-78;
sine[7351]=-78;
sine[7352]=-78;
sine[7353]=-78;
sine[7354]=-78;
sine[7355]=-78;
sine[7356]=-78;
sine[7357]=-78;
sine[7358]=-78;
sine[7359]=-78;
sine[7360]=-78;
sine[7361]=-78;
sine[7362]=-78;
sine[7363]=-78;
sine[7364]=-78;
sine[7365]=-78;
sine[7366]=-78;
sine[7367]=-78;
sine[7368]=-78;
sine[7369]=-78;
sine[7370]=-78;
sine[7371]=-78;
sine[7372]=-78;
sine[7373]=-78;
sine[7374]=-78;
sine[7375]=-78;
sine[7376]=-78;
sine[7377]=-78;
sine[7378]=-78;
sine[7379]=-78;
sine[7380]=-78;
sine[7381]=-78;
sine[7382]=-78;
sine[7383]=-78;
sine[7384]=-78;
sine[7385]=-78;
sine[7386]=-78;
sine[7387]=-78;
sine[7388]=-78;
sine[7389]=-78;
sine[7390]=-78;
sine[7391]=-78;
sine[7392]=-78;
sine[7393]=-78;
sine[7394]=-78;
sine[7395]=-78;
sine[7396]=-78;
sine[7397]=-78;
sine[7398]=-78;
sine[7399]=-78;
sine[7400]=-78;
sine[7401]=-78;
sine[7402]=-78;
sine[7403]=-78;
sine[7404]=-78;
sine[7405]=-78;
sine[7406]=-78;
sine[7407]=-78;
sine[7408]=-78;
sine[7409]=-78;
sine[7410]=-78;
sine[7411]=-78;
sine[7412]=-78;
sine[7413]=-78;
sine[7414]=-78;
sine[7415]=-78;
sine[7416]=-78;
sine[7417]=-78;
sine[7418]=-78;
sine[7419]=-78;
sine[7420]=-78;
sine[7421]=-78;
sine[7422]=-78;
sine[7423]=-78;
sine[7424]=-78;
sine[7425]=-78;
sine[7426]=-78;
sine[7427]=-78;
sine[7428]=-78;
sine[7429]=-78;
sine[7430]=-78;
sine[7431]=-78;
sine[7432]=-78;
sine[7433]=-78;
sine[7434]=-78;
sine[7435]=-78;
sine[7436]=-78;
sine[7437]=-78;
sine[7438]=-78;
sine[7439]=-78;
sine[7440]=-78;
sine[7441]=-78;
sine[7442]=-78;
sine[7443]=-78;
sine[7444]=-78;
sine[7445]=-78;
sine[7446]=-78;
sine[7447]=-78;
sine[7448]=-78;
sine[7449]=-78;
sine[7450]=-78;
sine[7451]=-78;
sine[7452]=-78;
sine[7453]=-78;
sine[7454]=-78;
sine[7455]=-78;
sine[7456]=-78;
sine[7457]=-78;
sine[7458]=-78;
sine[7459]=-78;
sine[7460]=-78;
sine[7461]=-78;
sine[7462]=-78;
sine[7463]=-78;
sine[7464]=-78;
sine[7465]=-78;
sine[7466]=-78;
sine[7467]=-78;
sine[7468]=-78;
sine[7469]=-78;
sine[7470]=-78;
sine[7471]=-78;
sine[7472]=-78;
sine[7473]=-78;
sine[7474]=-78;
sine[7475]=-78;
sine[7476]=-78;
sine[7477]=-78;
sine[7478]=-78;
sine[7479]=-78;
sine[7480]=-78;
sine[7481]=-78;
sine[7482]=-78;
sine[7483]=-78;
sine[7484]=-78;
sine[7485]=-78;
sine[7486]=-78;
sine[7487]=-78;
sine[7488]=-78;
sine[7489]=-78;
sine[7490]=-78;
sine[7491]=-78;
sine[7492]=-78;
sine[7493]=-78;
sine[7494]=-78;
sine[7495]=-78;
sine[7496]=-78;
sine[7497]=-78;
sine[7498]=-78;
sine[7499]=-78;
sine[7500]=-78;
sine[7501]=-78;
sine[7502]=-78;
sine[7503]=-78;
sine[7504]=-78;
sine[7505]=-78;
sine[7506]=-78;
sine[7507]=-78;
sine[7508]=-78;
sine[7509]=-78;
sine[7510]=-78;
sine[7511]=-78;
sine[7512]=-78;
sine[7513]=-78;
sine[7514]=-78;
sine[7515]=-78;
sine[7516]=-78;
sine[7517]=-78;
sine[7518]=-78;
sine[7519]=-78;
sine[7520]=-78;
sine[7521]=-78;
sine[7522]=-78;
sine[7523]=-78;
sine[7524]=-78;
sine[7525]=-78;
sine[7526]=-78;
sine[7527]=-78;
sine[7528]=-78;
sine[7529]=-78;
sine[7530]=-78;
sine[7531]=-78;
sine[7532]=-78;
sine[7533]=-78;
sine[7534]=-78;
sine[7535]=-78;
sine[7536]=-78;
sine[7537]=-78;
sine[7538]=-78;
sine[7539]=-78;
sine[7540]=-78;
sine[7541]=-78;
sine[7542]=-78;
sine[7543]=-78;
sine[7544]=-78;
sine[7545]=-78;
sine[7546]=-78;
sine[7547]=-78;
sine[7548]=-78;
sine[7549]=-78;
sine[7550]=-78;
sine[7551]=-78;
sine[7552]=-78;
sine[7553]=-78;
sine[7554]=-78;
sine[7555]=-78;
sine[7556]=-78;
sine[7557]=-78;
sine[7558]=-78;
sine[7559]=-78;
sine[7560]=-78;
sine[7561]=-78;
sine[7562]=-78;
sine[7563]=-78;
sine[7564]=-78;
sine[7565]=-78;
sine[7566]=-78;
sine[7567]=-78;
sine[7568]=-78;
sine[7569]=-78;
sine[7570]=-78;
sine[7571]=-78;
sine[7572]=-78;
sine[7573]=-78;
sine[7574]=-78;
sine[7575]=-78;
sine[7576]=-78;
sine[7577]=-78;
sine[7578]=-78;
sine[7579]=-78;
sine[7580]=-78;
sine[7581]=-78;
sine[7582]=-78;
sine[7583]=-78;
sine[7584]=-78;
sine[7585]=-78;
sine[7586]=-78;
sine[7587]=-78;
sine[7588]=-78;
sine[7589]=-78;
sine[7590]=-78;
sine[7591]=-78;
sine[7592]=-78;
sine[7593]=-78;
sine[7594]=-78;
sine[7595]=-78;
sine[7596]=-78;
sine[7597]=-78;
sine[7598]=-78;
sine[7599]=-78;
sine[7600]=-78;
sine[7601]=-78;
sine[7602]=-78;
sine[7603]=-78;
sine[7604]=-78;
sine[7605]=-78;
sine[7606]=-78;
sine[7607]=-78;
sine[7608]=-78;
sine[7609]=-78;
sine[7610]=-78;
sine[7611]=-78;
sine[7612]=-78;
sine[7613]=-78;
sine[7614]=-78;
sine[7615]=-78;
sine[7616]=-78;
sine[7617]=-78;
sine[7618]=-78;
sine[7619]=-78;
sine[7620]=-78;
sine[7621]=-78;
sine[7622]=-78;
sine[7623]=-78;
sine[7624]=-78;
sine[7625]=-78;
sine[7626]=-78;
sine[7627]=-78;
sine[7628]=-78;
sine[7629]=-78;
sine[7630]=-78;
sine[7631]=-78;
sine[7632]=-78;
sine[7633]=-78;
sine[7634]=-78;
sine[7635]=-78;
sine[7636]=-78;
sine[7637]=-78;
sine[7638]=-78;
sine[7639]=-78;
sine[7640]=-78;
sine[7641]=-78;
sine[7642]=-78;
sine[7643]=-78;
sine[7644]=-78;
sine[7645]=-78;
sine[7646]=-78;
sine[7647]=-78;
sine[7648]=-78;
sine[7649]=-78;
sine[7650]=-78;
sine[7651]=-78;
sine[7652]=-78;
sine[7653]=-78;
sine[7654]=-78;
sine[7655]=-78;
sine[7656]=-78;
sine[7657]=-78;
sine[7658]=-78;
sine[7659]=-78;
sine[7660]=-78;
sine[7661]=-78;
sine[7662]=-78;
sine[7663]=-78;
sine[7664]=-78;
sine[7665]=-78;
sine[7666]=-78;
sine[7667]=-78;
sine[7668]=-78;
sine[7669]=-78;
sine[7670]=-78;
sine[7671]=-78;
sine[7672]=-78;
sine[7673]=-78;
sine[7674]=-78;
sine[7675]=-78;
sine[7676]=-78;
sine[7677]=-78;
sine[7678]=-78;
sine[7679]=-78;
sine[7680]=-78;
sine[7681]=-78;
sine[7682]=-78;
sine[7683]=-78;
sine[7684]=-78;
sine[7685]=-78;
sine[7686]=-78;
sine[7687]=-78;
sine[7688]=-78;
sine[7689]=-78;
sine[7690]=-78;
sine[7691]=-78;
sine[7692]=-78;
sine[7693]=-78;
sine[7694]=-78;
sine[7695]=-78;
sine[7696]=-78;
sine[7697]=-78;
sine[7698]=-78;
sine[7699]=-78;
sine[7700]=-78;
sine[7701]=-78;
sine[7702]=-77;
sine[7703]=-77;
sine[7704]=-77;
sine[7705]=-77;
sine[7706]=-77;
sine[7707]=-77;
sine[7708]=-77;
sine[7709]=-77;
sine[7710]=-77;
sine[7711]=-77;
sine[7712]=-77;
sine[7713]=-77;
sine[7714]=-77;
sine[7715]=-77;
sine[7716]=-77;
sine[7717]=-77;
sine[7718]=-77;
sine[7719]=-77;
sine[7720]=-77;
sine[7721]=-77;
sine[7722]=-77;
sine[7723]=-77;
sine[7724]=-77;
sine[7725]=-77;
sine[7726]=-77;
sine[7727]=-77;
sine[7728]=-77;
sine[7729]=-77;
sine[7730]=-77;
sine[7731]=-77;
sine[7732]=-77;
sine[7733]=-77;
sine[7734]=-77;
sine[7735]=-77;
sine[7736]=-77;
sine[7737]=-77;
sine[7738]=-77;
sine[7739]=-77;
sine[7740]=-77;
sine[7741]=-77;
sine[7742]=-77;
sine[7743]=-77;
sine[7744]=-77;
sine[7745]=-77;
sine[7746]=-77;
sine[7747]=-77;
sine[7748]=-77;
sine[7749]=-77;
sine[7750]=-77;
sine[7751]=-77;
sine[7752]=-77;
sine[7753]=-77;
sine[7754]=-77;
sine[7755]=-77;
sine[7756]=-77;
sine[7757]=-77;
sine[7758]=-77;
sine[7759]=-77;
sine[7760]=-77;
sine[7761]=-77;
sine[7762]=-77;
sine[7763]=-77;
sine[7764]=-77;
sine[7765]=-77;
sine[7766]=-77;
sine[7767]=-77;
sine[7768]=-77;
sine[7769]=-77;
sine[7770]=-77;
sine[7771]=-77;
sine[7772]=-77;
sine[7773]=-77;
sine[7774]=-77;
sine[7775]=-77;
sine[7776]=-77;
sine[7777]=-77;
sine[7778]=-77;
sine[7779]=-77;
sine[7780]=-77;
sine[7781]=-77;
sine[7782]=-77;
sine[7783]=-77;
sine[7784]=-77;
sine[7785]=-77;
sine[7786]=-77;
sine[7787]=-77;
sine[7788]=-77;
sine[7789]=-77;
sine[7790]=-77;
sine[7791]=-77;
sine[7792]=-77;
sine[7793]=-77;
sine[7794]=-77;
sine[7795]=-77;
sine[7796]=-77;
sine[7797]=-77;
sine[7798]=-77;
sine[7799]=-77;
sine[7800]=-77;
sine[7801]=-77;
sine[7802]=-77;
sine[7803]=-77;
sine[7804]=-77;
sine[7805]=-77;
sine[7806]=-77;
sine[7807]=-77;
sine[7808]=-77;
sine[7809]=-77;
sine[7810]=-77;
sine[7811]=-77;
sine[7812]=-77;
sine[7813]=-77;
sine[7814]=-77;
sine[7815]=-77;
sine[7816]=-77;
sine[7817]=-77;
sine[7818]=-77;
sine[7819]=-77;
sine[7820]=-77;
sine[7821]=-77;
sine[7822]=-77;
sine[7823]=-77;
sine[7824]=-77;
sine[7825]=-77;
sine[7826]=-76;
sine[7827]=-76;
sine[7828]=-76;
sine[7829]=-76;
sine[7830]=-76;
sine[7831]=-76;
sine[7832]=-76;
sine[7833]=-76;
sine[7834]=-76;
sine[7835]=-76;
sine[7836]=-76;
sine[7837]=-76;
sine[7838]=-76;
sine[7839]=-76;
sine[7840]=-76;
sine[7841]=-76;
sine[7842]=-76;
sine[7843]=-76;
sine[7844]=-76;
sine[7845]=-76;
sine[7846]=-76;
sine[7847]=-76;
sine[7848]=-76;
sine[7849]=-76;
sine[7850]=-76;
sine[7851]=-76;
sine[7852]=-76;
sine[7853]=-76;
sine[7854]=-76;
sine[7855]=-76;
sine[7856]=-76;
sine[7857]=-76;
sine[7858]=-76;
sine[7859]=-76;
sine[7860]=-76;
sine[7861]=-76;
sine[7862]=-76;
sine[7863]=-76;
sine[7864]=-76;
sine[7865]=-76;
sine[7866]=-76;
sine[7867]=-76;
sine[7868]=-76;
sine[7869]=-76;
sine[7870]=-76;
sine[7871]=-76;
sine[7872]=-76;
sine[7873]=-76;
sine[7874]=-76;
sine[7875]=-76;
sine[7876]=-76;
sine[7877]=-76;
sine[7878]=-76;
sine[7879]=-76;
sine[7880]=-76;
sine[7881]=-76;
sine[7882]=-76;
sine[7883]=-76;
sine[7884]=-76;
sine[7885]=-76;
sine[7886]=-76;
sine[7887]=-76;
sine[7888]=-76;
sine[7889]=-76;
sine[7890]=-76;
sine[7891]=-76;
sine[7892]=-76;
sine[7893]=-76;
sine[7894]=-76;
sine[7895]=-76;
sine[7896]=-76;
sine[7897]=-76;
sine[7898]=-76;
sine[7899]=-76;
sine[7900]=-76;
sine[7901]=-76;
sine[7902]=-76;
sine[7903]=-76;
sine[7904]=-76;
sine[7905]=-76;
sine[7906]=-76;
sine[7907]=-76;
sine[7908]=-76;
sine[7909]=-76;
sine[7910]=-76;
sine[7911]=-76;
sine[7912]=-76;
sine[7913]=-76;
sine[7914]=-75;
sine[7915]=-75;
sine[7916]=-75;
sine[7917]=-75;
sine[7918]=-75;
sine[7919]=-75;
sine[7920]=-75;
sine[7921]=-75;
sine[7922]=-75;
sine[7923]=-75;
sine[7924]=-75;
sine[7925]=-75;
sine[7926]=-75;
sine[7927]=-75;
sine[7928]=-75;
sine[7929]=-75;
sine[7930]=-75;
sine[7931]=-75;
sine[7932]=-75;
sine[7933]=-75;
sine[7934]=-75;
sine[7935]=-75;
sine[7936]=-75;
sine[7937]=-75;
sine[7938]=-75;
sine[7939]=-75;
sine[7940]=-75;
sine[7941]=-75;
sine[7942]=-75;
sine[7943]=-75;
sine[7944]=-75;
sine[7945]=-75;
sine[7946]=-75;
sine[7947]=-75;
sine[7948]=-75;
sine[7949]=-75;
sine[7950]=-75;
sine[7951]=-75;
sine[7952]=-75;
sine[7953]=-75;
sine[7954]=-75;
sine[7955]=-75;
sine[7956]=-75;
sine[7957]=-75;
sine[7958]=-75;
sine[7959]=-75;
sine[7960]=-75;
sine[7961]=-75;
sine[7962]=-75;
sine[7963]=-75;
sine[7964]=-75;
sine[7965]=-75;
sine[7966]=-75;
sine[7967]=-75;
sine[7968]=-75;
sine[7969]=-75;
sine[7970]=-75;
sine[7971]=-75;
sine[7972]=-75;
sine[7973]=-75;
sine[7974]=-75;
sine[7975]=-75;
sine[7976]=-75;
sine[7977]=-75;
sine[7978]=-75;
sine[7979]=-75;
sine[7980]=-75;
sine[7981]=-75;
sine[7982]=-75;
sine[7983]=-75;
sine[7984]=-75;
sine[7985]=-75;
sine[7986]=-75;
sine[7987]=-74;
sine[7988]=-74;
sine[7989]=-74;
sine[7990]=-74;
sine[7991]=-74;
sine[7992]=-74;
sine[7993]=-74;
sine[7994]=-74;
sine[7995]=-74;
sine[7996]=-74;
sine[7997]=-74;
sine[7998]=-74;
sine[7999]=-74;
sine[8000]=-74;
sine[8001]=-74;
sine[8002]=-74;
sine[8003]=-74;
sine[8004]=-74;
sine[8005]=-74;
sine[8006]=-74;
sine[8007]=-74;
sine[8008]=-74;
sine[8009]=-74;
sine[8010]=-74;
sine[8011]=-74;
sine[8012]=-74;
sine[8013]=-74;
sine[8014]=-74;
sine[8015]=-74;
sine[8016]=-74;
sine[8017]=-74;
sine[8018]=-74;
sine[8019]=-74;
sine[8020]=-74;
sine[8021]=-74;
sine[8022]=-74;
sine[8023]=-74;
sine[8024]=-74;
sine[8025]=-74;
sine[8026]=-74;
sine[8027]=-74;
sine[8028]=-74;
sine[8029]=-74;
sine[8030]=-74;
sine[8031]=-74;
sine[8032]=-74;
sine[8033]=-74;
sine[8034]=-74;
sine[8035]=-74;
sine[8036]=-74;
sine[8037]=-74;
sine[8038]=-74;
sine[8039]=-74;
sine[8040]=-74;
sine[8041]=-74;
sine[8042]=-74;
sine[8043]=-74;
sine[8044]=-74;
sine[8045]=-74;
sine[8046]=-74;
sine[8047]=-74;
sine[8048]=-74;
sine[8049]=-74;
sine[8050]=-74;
sine[8051]=-73;
sine[8052]=-73;
sine[8053]=-73;
sine[8054]=-73;
sine[8055]=-73;
sine[8056]=-73;
sine[8057]=-73;
sine[8058]=-73;
sine[8059]=-73;
sine[8060]=-73;
sine[8061]=-73;
sine[8062]=-73;
sine[8063]=-73;
sine[8064]=-73;
sine[8065]=-73;
sine[8066]=-73;
sine[8067]=-73;
sine[8068]=-73;
sine[8069]=-73;
sine[8070]=-73;
sine[8071]=-73;
sine[8072]=-73;
sine[8073]=-73;
sine[8074]=-73;
sine[8075]=-73;
sine[8076]=-73;
sine[8077]=-73;
sine[8078]=-73;
sine[8079]=-73;
sine[8080]=-73;
sine[8081]=-73;
sine[8082]=-73;
sine[8083]=-73;
sine[8084]=-73;
sine[8085]=-73;
sine[8086]=-73;
sine[8087]=-73;
sine[8088]=-73;
sine[8089]=-73;
sine[8090]=-73;
sine[8091]=-73;
sine[8092]=-73;
sine[8093]=-73;
sine[8094]=-73;
sine[8095]=-73;
sine[8096]=-73;
sine[8097]=-73;
sine[8098]=-73;
sine[8099]=-73;
sine[8100]=-73;
sine[8101]=-73;
sine[8102]=-73;
sine[8103]=-73;
sine[8104]=-73;
sine[8105]=-73;
sine[8106]=-73;
sine[8107]=-73;
sine[8108]=-72;
sine[8109]=-72;
sine[8110]=-72;
sine[8111]=-72;
sine[8112]=-72;
sine[8113]=-72;
sine[8114]=-72;
sine[8115]=-72;
sine[8116]=-72;
sine[8117]=-72;
sine[8118]=-72;
sine[8119]=-72;
sine[8120]=-72;
sine[8121]=-72;
sine[8122]=-72;
sine[8123]=-72;
sine[8124]=-72;
sine[8125]=-72;
sine[8126]=-72;
sine[8127]=-72;
sine[8128]=-72;
sine[8129]=-72;
sine[8130]=-72;
sine[8131]=-72;
sine[8132]=-72;
sine[8133]=-72;
sine[8134]=-72;
sine[8135]=-72;
sine[8136]=-72;
sine[8137]=-72;
sine[8138]=-72;
sine[8139]=-72;
sine[8140]=-72;
sine[8141]=-72;
sine[8142]=-72;
sine[8143]=-72;
sine[8144]=-72;
sine[8145]=-72;
sine[8146]=-72;
sine[8147]=-72;
sine[8148]=-72;
sine[8149]=-72;
sine[8150]=-72;
sine[8151]=-72;
sine[8152]=-72;
sine[8153]=-72;
sine[8154]=-72;
sine[8155]=-72;
sine[8156]=-72;
sine[8157]=-72;
sine[8158]=-72;
sine[8159]=-72;
sine[8160]=-72;
sine[8161]=-71;
sine[8162]=-71;
sine[8163]=-71;
sine[8164]=-71;
sine[8165]=-71;
sine[8166]=-71;
sine[8167]=-71;
sine[8168]=-71;
sine[8169]=-71;
sine[8170]=-71;
sine[8171]=-71;
sine[8172]=-71;
sine[8173]=-71;
sine[8174]=-71;
sine[8175]=-71;
sine[8176]=-71;
sine[8177]=-71;
sine[8178]=-71;
sine[8179]=-71;
sine[8180]=-71;
sine[8181]=-71;
sine[8182]=-71;
sine[8183]=-71;
sine[8184]=-71;
sine[8185]=-71;
sine[8186]=-71;
sine[8187]=-71;
sine[8188]=-71;
sine[8189]=-71;
sine[8190]=-71;
sine[8191]=-71;
sine[8192]=-71;
sine[8193]=-71;
sine[8194]=-71;
sine[8195]=-71;
sine[8196]=-71;
sine[8197]=-71;
sine[8198]=-71;
sine[8199]=-71;
sine[8200]=-71;
sine[8201]=-71;
sine[8202]=-71;
sine[8203]=-71;
sine[8204]=-71;
sine[8205]=-71;
sine[8206]=-71;
sine[8207]=-71;
sine[8208]=-71;
sine[8209]=-71;
sine[8210]=-70;
sine[8211]=-70;
sine[8212]=-70;
sine[8213]=-70;
sine[8214]=-70;
sine[8215]=-70;
sine[8216]=-70;
sine[8217]=-70;
sine[8218]=-70;
sine[8219]=-70;
sine[8220]=-70;
sine[8221]=-70;
sine[8222]=-70;
sine[8223]=-70;
sine[8224]=-70;
sine[8225]=-70;
sine[8226]=-70;
sine[8227]=-70;
sine[8228]=-70;
sine[8229]=-70;
sine[8230]=-70;
sine[8231]=-70;
sine[8232]=-70;
sine[8233]=-70;
sine[8234]=-70;
sine[8235]=-70;
sine[8236]=-70;
sine[8237]=-70;
sine[8238]=-70;
sine[8239]=-70;
sine[8240]=-70;
sine[8241]=-70;
sine[8242]=-70;
sine[8243]=-70;
sine[8244]=-70;
sine[8245]=-70;
sine[8246]=-70;
sine[8247]=-70;
sine[8248]=-70;
sine[8249]=-70;
sine[8250]=-70;
sine[8251]=-70;
sine[8252]=-70;
sine[8253]=-70;
sine[8254]=-70;
sine[8255]=-69;
sine[8256]=-69;
sine[8257]=-69;
sine[8258]=-69;
sine[8259]=-69;
sine[8260]=-69;
sine[8261]=-69;
sine[8262]=-69;
sine[8263]=-69;
sine[8264]=-69;
sine[8265]=-69;
sine[8266]=-69;
sine[8267]=-69;
sine[8268]=-69;
sine[8269]=-69;
sine[8270]=-69;
sine[8271]=-69;
sine[8272]=-69;
sine[8273]=-69;
sine[8274]=-69;
sine[8275]=-69;
sine[8276]=-69;
sine[8277]=-69;
sine[8278]=-69;
sine[8279]=-69;
sine[8280]=-69;
sine[8281]=-69;
sine[8282]=-69;
sine[8283]=-69;
sine[8284]=-69;
sine[8285]=-69;
sine[8286]=-69;
sine[8287]=-69;
sine[8288]=-69;
sine[8289]=-69;
sine[8290]=-69;
sine[8291]=-69;
sine[8292]=-69;
sine[8293]=-69;
sine[8294]=-69;
sine[8295]=-69;
sine[8296]=-69;
sine[8297]=-69;
sine[8298]=-69;
sine[8299]=-68;
sine[8300]=-68;
sine[8301]=-68;
sine[8302]=-68;
sine[8303]=-68;
sine[8304]=-68;
sine[8305]=-68;
sine[8306]=-68;
sine[8307]=-68;
sine[8308]=-68;
sine[8309]=-68;
sine[8310]=-68;
sine[8311]=-68;
sine[8312]=-68;
sine[8313]=-68;
sine[8314]=-68;
sine[8315]=-68;
sine[8316]=-68;
sine[8317]=-68;
sine[8318]=-68;
sine[8319]=-68;
sine[8320]=-68;
sine[8321]=-68;
sine[8322]=-68;
sine[8323]=-68;
sine[8324]=-68;
sine[8325]=-68;
sine[8326]=-68;
sine[8327]=-68;
sine[8328]=-68;
sine[8329]=-68;
sine[8330]=-68;
sine[8331]=-68;
sine[8332]=-68;
sine[8333]=-68;
sine[8334]=-68;
sine[8335]=-68;
sine[8336]=-68;
sine[8337]=-68;
sine[8338]=-68;
sine[8339]=-68;
sine[8340]=-67;
sine[8341]=-67;
sine[8342]=-67;
sine[8343]=-67;
sine[8344]=-67;
sine[8345]=-67;
sine[8346]=-67;
sine[8347]=-67;
sine[8348]=-67;
sine[8349]=-67;
sine[8350]=-67;
sine[8351]=-67;
sine[8352]=-67;
sine[8353]=-67;
sine[8354]=-67;
sine[8355]=-67;
sine[8356]=-67;
sine[8357]=-67;
sine[8358]=-67;
sine[8359]=-67;
sine[8360]=-67;
sine[8361]=-67;
sine[8362]=-67;
sine[8363]=-67;
sine[8364]=-67;
sine[8365]=-67;
sine[8366]=-67;
sine[8367]=-67;
sine[8368]=-67;
sine[8369]=-67;
sine[8370]=-67;
sine[8371]=-67;
sine[8372]=-67;
sine[8373]=-67;
sine[8374]=-67;
sine[8375]=-67;
sine[8376]=-67;
sine[8377]=-67;
sine[8378]=-67;
sine[8379]=-67;
sine[8380]=-66;
sine[8381]=-66;
sine[8382]=-66;
sine[8383]=-66;
sine[8384]=-66;
sine[8385]=-66;
sine[8386]=-66;
sine[8387]=-66;
sine[8388]=-66;
sine[8389]=-66;
sine[8390]=-66;
sine[8391]=-66;
sine[8392]=-66;
sine[8393]=-66;
sine[8394]=-66;
sine[8395]=-66;
sine[8396]=-66;
sine[8397]=-66;
sine[8398]=-66;
sine[8399]=-66;
sine[8400]=-66;
sine[8401]=-66;
sine[8402]=-66;
sine[8403]=-66;
sine[8404]=-66;
sine[8405]=-66;
sine[8406]=-66;
sine[8407]=-66;
sine[8408]=-66;
sine[8409]=-66;
sine[8410]=-66;
sine[8411]=-66;
sine[8412]=-66;
sine[8413]=-66;
sine[8414]=-66;
sine[8415]=-66;
sine[8416]=-66;
sine[8417]=-66;
sine[8418]=-65;
sine[8419]=-65;
sine[8420]=-65;
sine[8421]=-65;
sine[8422]=-65;
sine[8423]=-65;
sine[8424]=-65;
sine[8425]=-65;
sine[8426]=-65;
sine[8427]=-65;
sine[8428]=-65;
sine[8429]=-65;
sine[8430]=-65;
sine[8431]=-65;
sine[8432]=-65;
sine[8433]=-65;
sine[8434]=-65;
sine[8435]=-65;
sine[8436]=-65;
sine[8437]=-65;
sine[8438]=-65;
sine[8439]=-65;
sine[8440]=-65;
sine[8441]=-65;
sine[8442]=-65;
sine[8443]=-65;
sine[8444]=-65;
sine[8445]=-65;
sine[8446]=-65;
sine[8447]=-65;
sine[8448]=-65;
sine[8449]=-65;
sine[8450]=-65;
sine[8451]=-65;
sine[8452]=-65;
sine[8453]=-65;
sine[8454]=-65;
sine[8455]=-64;
sine[8456]=-64;
sine[8457]=-64;
sine[8458]=-64;
sine[8459]=-64;
sine[8460]=-64;
sine[8461]=-64;
sine[8462]=-64;
sine[8463]=-64;
sine[8464]=-64;
sine[8465]=-64;
sine[8466]=-64;
sine[8467]=-64;
sine[8468]=-64;
sine[8469]=-64;
sine[8470]=-64;
sine[8471]=-64;
sine[8472]=-64;
sine[8473]=-64;
sine[8474]=-64;
sine[8475]=-64;
sine[8476]=-64;
sine[8477]=-64;
sine[8478]=-64;
sine[8479]=-64;
sine[8480]=-64;
sine[8481]=-64;
sine[8482]=-64;
sine[8483]=-64;
sine[8484]=-64;
sine[8485]=-64;
sine[8486]=-64;
sine[8487]=-64;
sine[8488]=-64;
sine[8489]=-64;
sine[8490]=-63;
sine[8491]=-63;
sine[8492]=-63;
sine[8493]=-63;
sine[8494]=-63;
sine[8495]=-63;
sine[8496]=-63;
sine[8497]=-63;
sine[8498]=-63;
sine[8499]=-63;
sine[8500]=-63;
sine[8501]=-63;
sine[8502]=-63;
sine[8503]=-63;
sine[8504]=-63;
sine[8505]=-63;
sine[8506]=-63;
sine[8507]=-63;
sine[8508]=-63;
sine[8509]=-63;
sine[8510]=-63;
sine[8511]=-63;
sine[8512]=-63;
sine[8513]=-63;
sine[8514]=-63;
sine[8515]=-63;
sine[8516]=-63;
sine[8517]=-63;
sine[8518]=-63;
sine[8519]=-63;
sine[8520]=-63;
sine[8521]=-63;
sine[8522]=-63;
sine[8523]=-63;
sine[8524]=-63;
sine[8525]=-62;
sine[8526]=-62;
sine[8527]=-62;
sine[8528]=-62;
sine[8529]=-62;
sine[8530]=-62;
sine[8531]=-62;
sine[8532]=-62;
sine[8533]=-62;
sine[8534]=-62;
sine[8535]=-62;
sine[8536]=-62;
sine[8537]=-62;
sine[8538]=-62;
sine[8539]=-62;
sine[8540]=-62;
sine[8541]=-62;
sine[8542]=-62;
sine[8543]=-62;
sine[8544]=-62;
sine[8545]=-62;
sine[8546]=-62;
sine[8547]=-62;
sine[8548]=-62;
sine[8549]=-62;
sine[8550]=-62;
sine[8551]=-62;
sine[8552]=-62;
sine[8553]=-62;
sine[8554]=-62;
sine[8555]=-62;
sine[8556]=-62;
sine[8557]=-62;
sine[8558]=-61;
sine[8559]=-61;
sine[8560]=-61;
sine[8561]=-61;
sine[8562]=-61;
sine[8563]=-61;
sine[8564]=-61;
sine[8565]=-61;
sine[8566]=-61;
sine[8567]=-61;
sine[8568]=-61;
sine[8569]=-61;
sine[8570]=-61;
sine[8571]=-61;
sine[8572]=-61;
sine[8573]=-61;
sine[8574]=-61;
sine[8575]=-61;
sine[8576]=-61;
sine[8577]=-61;
sine[8578]=-61;
sine[8579]=-61;
sine[8580]=-61;
sine[8581]=-61;
sine[8582]=-61;
sine[8583]=-61;
sine[8584]=-61;
sine[8585]=-61;
sine[8586]=-61;
sine[8587]=-61;
sine[8588]=-61;
sine[8589]=-61;
sine[8590]=-61;
sine[8591]=-60;
sine[8592]=-60;
sine[8593]=-60;
sine[8594]=-60;
sine[8595]=-60;
sine[8596]=-60;
sine[8597]=-60;
sine[8598]=-60;
sine[8599]=-60;
sine[8600]=-60;
sine[8601]=-60;
sine[8602]=-60;
sine[8603]=-60;
sine[8604]=-60;
sine[8605]=-60;
sine[8606]=-60;
sine[8607]=-60;
sine[8608]=-60;
sine[8609]=-60;
sine[8610]=-60;
sine[8611]=-60;
sine[8612]=-60;
sine[8613]=-60;
sine[8614]=-60;
sine[8615]=-60;
sine[8616]=-60;
sine[8617]=-60;
sine[8618]=-60;
sine[8619]=-60;
sine[8620]=-60;
sine[8621]=-60;
sine[8622]=-60;
sine[8623]=-59;
sine[8624]=-59;
sine[8625]=-59;
sine[8626]=-59;
sine[8627]=-59;
sine[8628]=-59;
sine[8629]=-59;
sine[8630]=-59;
sine[8631]=-59;
sine[8632]=-59;
sine[8633]=-59;
sine[8634]=-59;
sine[8635]=-59;
sine[8636]=-59;
sine[8637]=-59;
sine[8638]=-59;
sine[8639]=-59;
sine[8640]=-59;
sine[8641]=-59;
sine[8642]=-59;
sine[8643]=-59;
sine[8644]=-59;
sine[8645]=-59;
sine[8646]=-59;
sine[8647]=-59;
sine[8648]=-59;
sine[8649]=-59;
sine[8650]=-59;
sine[8651]=-59;
sine[8652]=-59;
sine[8653]=-59;
sine[8654]=-58;
sine[8655]=-58;
sine[8656]=-58;
sine[8657]=-58;
sine[8658]=-58;
sine[8659]=-58;
sine[8660]=-58;
sine[8661]=-58;
sine[8662]=-58;
sine[8663]=-58;
sine[8664]=-58;
sine[8665]=-58;
sine[8666]=-58;
sine[8667]=-58;
sine[8668]=-58;
sine[8669]=-58;
sine[8670]=-58;
sine[8671]=-58;
sine[8672]=-58;
sine[8673]=-58;
sine[8674]=-58;
sine[8675]=-58;
sine[8676]=-58;
sine[8677]=-58;
sine[8678]=-58;
sine[8679]=-58;
sine[8680]=-58;
sine[8681]=-58;
sine[8682]=-58;
sine[8683]=-58;
sine[8684]=-57;
sine[8685]=-57;
sine[8686]=-57;
sine[8687]=-57;
sine[8688]=-57;
sine[8689]=-57;
sine[8690]=-57;
sine[8691]=-57;
sine[8692]=-57;
sine[8693]=-57;
sine[8694]=-57;
sine[8695]=-57;
sine[8696]=-57;
sine[8697]=-57;
sine[8698]=-57;
sine[8699]=-57;
sine[8700]=-57;
sine[8701]=-57;
sine[8702]=-57;
sine[8703]=-57;
sine[8704]=-57;
sine[8705]=-57;
sine[8706]=-57;
sine[8707]=-57;
sine[8708]=-57;
sine[8709]=-57;
sine[8710]=-57;
sine[8711]=-57;
sine[8712]=-57;
sine[8713]=-57;
sine[8714]=-56;
sine[8715]=-56;
sine[8716]=-56;
sine[8717]=-56;
sine[8718]=-56;
sine[8719]=-56;
sine[8720]=-56;
sine[8721]=-56;
sine[8722]=-56;
sine[8723]=-56;
sine[8724]=-56;
sine[8725]=-56;
sine[8726]=-56;
sine[8727]=-56;
sine[8728]=-56;
sine[8729]=-56;
sine[8730]=-56;
sine[8731]=-56;
sine[8732]=-56;
sine[8733]=-56;
sine[8734]=-56;
sine[8735]=-56;
sine[8736]=-56;
sine[8737]=-56;
sine[8738]=-56;
sine[8739]=-56;
sine[8740]=-56;
sine[8741]=-56;
sine[8742]=-56;
sine[8743]=-55;
sine[8744]=-55;
sine[8745]=-55;
sine[8746]=-55;
sine[8747]=-55;
sine[8748]=-55;
sine[8749]=-55;
sine[8750]=-55;
sine[8751]=-55;
sine[8752]=-55;
sine[8753]=-55;
sine[8754]=-55;
sine[8755]=-55;
sine[8756]=-55;
sine[8757]=-55;
sine[8758]=-55;
sine[8759]=-55;
sine[8760]=-55;
sine[8761]=-55;
sine[8762]=-55;
sine[8763]=-55;
sine[8764]=-55;
sine[8765]=-55;
sine[8766]=-55;
sine[8767]=-55;
sine[8768]=-55;
sine[8769]=-55;
sine[8770]=-55;
sine[8771]=-55;
sine[8772]=-54;
sine[8773]=-54;
sine[8774]=-54;
sine[8775]=-54;
sine[8776]=-54;
sine[8777]=-54;
sine[8778]=-54;
sine[8779]=-54;
sine[8780]=-54;
sine[8781]=-54;
sine[8782]=-54;
sine[8783]=-54;
sine[8784]=-54;
sine[8785]=-54;
sine[8786]=-54;
sine[8787]=-54;
sine[8788]=-54;
sine[8789]=-54;
sine[8790]=-54;
sine[8791]=-54;
sine[8792]=-54;
sine[8793]=-54;
sine[8794]=-54;
sine[8795]=-54;
sine[8796]=-54;
sine[8797]=-54;
sine[8798]=-54;
sine[8799]=-54;
sine[8800]=-53;
sine[8801]=-53;
sine[8802]=-53;
sine[8803]=-53;
sine[8804]=-53;
sine[8805]=-53;
sine[8806]=-53;
sine[8807]=-53;
sine[8808]=-53;
sine[8809]=-53;
sine[8810]=-53;
sine[8811]=-53;
sine[8812]=-53;
sine[8813]=-53;
sine[8814]=-53;
sine[8815]=-53;
sine[8816]=-53;
sine[8817]=-53;
sine[8818]=-53;
sine[8819]=-53;
sine[8820]=-53;
sine[8821]=-53;
sine[8822]=-53;
sine[8823]=-53;
sine[8824]=-53;
sine[8825]=-53;
sine[8826]=-53;
sine[8827]=-53;
sine[8828]=-52;
sine[8829]=-52;
sine[8830]=-52;
sine[8831]=-52;
sine[8832]=-52;
sine[8833]=-52;
sine[8834]=-52;
sine[8835]=-52;
sine[8836]=-52;
sine[8837]=-52;
sine[8838]=-52;
sine[8839]=-52;
sine[8840]=-52;
sine[8841]=-52;
sine[8842]=-52;
sine[8843]=-52;
sine[8844]=-52;
sine[8845]=-52;
sine[8846]=-52;
sine[8847]=-52;
sine[8848]=-52;
sine[8849]=-52;
sine[8850]=-52;
sine[8851]=-52;
sine[8852]=-52;
sine[8853]=-52;
sine[8854]=-52;
sine[8855]=-51;
sine[8856]=-51;
sine[8857]=-51;
sine[8858]=-51;
sine[8859]=-51;
sine[8860]=-51;
sine[8861]=-51;
sine[8862]=-51;
sine[8863]=-51;
sine[8864]=-51;
sine[8865]=-51;
sine[8866]=-51;
sine[8867]=-51;
sine[8868]=-51;
sine[8869]=-51;
sine[8870]=-51;
sine[8871]=-51;
sine[8872]=-51;
sine[8873]=-51;
sine[8874]=-51;
sine[8875]=-51;
sine[8876]=-51;
sine[8877]=-51;
sine[8878]=-51;
sine[8879]=-51;
sine[8880]=-51;
sine[8881]=-51;
sine[8882]=-50;
sine[8883]=-50;
sine[8884]=-50;
sine[8885]=-50;
sine[8886]=-50;
sine[8887]=-50;
sine[8888]=-50;
sine[8889]=-50;
sine[8890]=-50;
sine[8891]=-50;
sine[8892]=-50;
sine[8893]=-50;
sine[8894]=-50;
sine[8895]=-50;
sine[8896]=-50;
sine[8897]=-50;
sine[8898]=-50;
sine[8899]=-50;
sine[8900]=-50;
sine[8901]=-50;
sine[8902]=-50;
sine[8903]=-50;
sine[8904]=-50;
sine[8905]=-50;
sine[8906]=-50;
sine[8907]=-50;
sine[8908]=-49;
sine[8909]=-49;
sine[8910]=-49;
sine[8911]=-49;
sine[8912]=-49;
sine[8913]=-49;
sine[8914]=-49;
sine[8915]=-49;
sine[8916]=-49;
sine[8917]=-49;
sine[8918]=-49;
sine[8919]=-49;
sine[8920]=-49;
sine[8921]=-49;
sine[8922]=-49;
sine[8923]=-49;
sine[8924]=-49;
sine[8925]=-49;
sine[8926]=-49;
sine[8927]=-49;
sine[8928]=-49;
sine[8929]=-49;
sine[8930]=-49;
sine[8931]=-49;
sine[8932]=-49;
sine[8933]=-49;
sine[8934]=-49;
sine[8935]=-48;
sine[8936]=-48;
sine[8937]=-48;
sine[8938]=-48;
sine[8939]=-48;
sine[8940]=-48;
sine[8941]=-48;
sine[8942]=-48;
sine[8943]=-48;
sine[8944]=-48;
sine[8945]=-48;
sine[8946]=-48;
sine[8947]=-48;
sine[8948]=-48;
sine[8949]=-48;
sine[8950]=-48;
sine[8951]=-48;
sine[8952]=-48;
sine[8953]=-48;
sine[8954]=-48;
sine[8955]=-48;
sine[8956]=-48;
sine[8957]=-48;
sine[8958]=-48;
sine[8959]=-48;
sine[8960]=-47;
sine[8961]=-47;
sine[8962]=-47;
sine[8963]=-47;
sine[8964]=-47;
sine[8965]=-47;
sine[8966]=-47;
sine[8967]=-47;
sine[8968]=-47;
sine[8969]=-47;
sine[8970]=-47;
sine[8971]=-47;
sine[8972]=-47;
sine[8973]=-47;
sine[8974]=-47;
sine[8975]=-47;
sine[8976]=-47;
sine[8977]=-47;
sine[8978]=-47;
sine[8979]=-47;
sine[8980]=-47;
sine[8981]=-47;
sine[8982]=-47;
sine[8983]=-47;
sine[8984]=-47;
sine[8985]=-47;
sine[8986]=-46;
sine[8987]=-46;
sine[8988]=-46;
sine[8989]=-46;
sine[8990]=-46;
sine[8991]=-46;
sine[8992]=-46;
sine[8993]=-46;
sine[8994]=-46;
sine[8995]=-46;
sine[8996]=-46;
sine[8997]=-46;
sine[8998]=-46;
sine[8999]=-46;
sine[9000]=-46;
sine[9001]=-46;
sine[9002]=-46;
sine[9003]=-46;
sine[9004]=-46;
sine[9005]=-46;
sine[9006]=-46;
sine[9007]=-46;
sine[9008]=-46;
sine[9009]=-46;
sine[9010]=-46;
sine[9011]=-45;
sine[9012]=-45;
sine[9013]=-45;
sine[9014]=-45;
sine[9015]=-45;
sine[9016]=-45;
sine[9017]=-45;
sine[9018]=-45;
sine[9019]=-45;
sine[9020]=-45;
sine[9021]=-45;
sine[9022]=-45;
sine[9023]=-45;
sine[9024]=-45;
sine[9025]=-45;
sine[9026]=-45;
sine[9027]=-45;
sine[9028]=-45;
sine[9029]=-45;
sine[9030]=-45;
sine[9031]=-45;
sine[9032]=-45;
sine[9033]=-45;
sine[9034]=-45;
sine[9035]=-45;
sine[9036]=-44;
sine[9037]=-44;
sine[9038]=-44;
sine[9039]=-44;
sine[9040]=-44;
sine[9041]=-44;
sine[9042]=-44;
sine[9043]=-44;
sine[9044]=-44;
sine[9045]=-44;
sine[9046]=-44;
sine[9047]=-44;
sine[9048]=-44;
sine[9049]=-44;
sine[9050]=-44;
sine[9051]=-44;
sine[9052]=-44;
sine[9053]=-44;
sine[9054]=-44;
sine[9055]=-44;
sine[9056]=-44;
sine[9057]=-44;
sine[9058]=-44;
sine[9059]=-44;
sine[9060]=-44;
sine[9061]=-43;
sine[9062]=-43;
sine[9063]=-43;
sine[9064]=-43;
sine[9065]=-43;
sine[9066]=-43;
sine[9067]=-43;
sine[9068]=-43;
sine[9069]=-43;
sine[9070]=-43;
sine[9071]=-43;
sine[9072]=-43;
sine[9073]=-43;
sine[9074]=-43;
sine[9075]=-43;
sine[9076]=-43;
sine[9077]=-43;
sine[9078]=-43;
sine[9079]=-43;
sine[9080]=-43;
sine[9081]=-43;
sine[9082]=-43;
sine[9083]=-43;
sine[9084]=-43;
sine[9085]=-42;
sine[9086]=-42;
sine[9087]=-42;
sine[9088]=-42;
sine[9089]=-42;
sine[9090]=-42;
sine[9091]=-42;
sine[9092]=-42;
sine[9093]=-42;
sine[9094]=-42;
sine[9095]=-42;
sine[9096]=-42;
sine[9097]=-42;
sine[9098]=-42;
sine[9099]=-42;
sine[9100]=-42;
sine[9101]=-42;
sine[9102]=-42;
sine[9103]=-42;
sine[9104]=-42;
sine[9105]=-42;
sine[9106]=-42;
sine[9107]=-42;
sine[9108]=-42;
sine[9109]=-41;
sine[9110]=-41;
sine[9111]=-41;
sine[9112]=-41;
sine[9113]=-41;
sine[9114]=-41;
sine[9115]=-41;
sine[9116]=-41;
sine[9117]=-41;
sine[9118]=-41;
sine[9119]=-41;
sine[9120]=-41;
sine[9121]=-41;
sine[9122]=-41;
sine[9123]=-41;
sine[9124]=-41;
sine[9125]=-41;
sine[9126]=-41;
sine[9127]=-41;
sine[9128]=-41;
sine[9129]=-41;
sine[9130]=-41;
sine[9131]=-41;
sine[9132]=-41;
sine[9133]=-40;
sine[9134]=-40;
sine[9135]=-40;
sine[9136]=-40;
sine[9137]=-40;
sine[9138]=-40;
sine[9139]=-40;
sine[9140]=-40;
sine[9141]=-40;
sine[9142]=-40;
sine[9143]=-40;
sine[9144]=-40;
sine[9145]=-40;
sine[9146]=-40;
sine[9147]=-40;
sine[9148]=-40;
sine[9149]=-40;
sine[9150]=-40;
sine[9151]=-40;
sine[9152]=-40;
sine[9153]=-40;
sine[9154]=-40;
sine[9155]=-40;
sine[9156]=-40;
sine[9157]=-39;
sine[9158]=-39;
sine[9159]=-39;
sine[9160]=-39;
sine[9161]=-39;
sine[9162]=-39;
sine[9163]=-39;
sine[9164]=-39;
sine[9165]=-39;
sine[9166]=-39;
sine[9167]=-39;
sine[9168]=-39;
sine[9169]=-39;
sine[9170]=-39;
sine[9171]=-39;
sine[9172]=-39;
sine[9173]=-39;
sine[9174]=-39;
sine[9175]=-39;
sine[9176]=-39;
sine[9177]=-39;
sine[9178]=-39;
sine[9179]=-39;
sine[9180]=-38;
sine[9181]=-38;
sine[9182]=-38;
sine[9183]=-38;
sine[9184]=-38;
sine[9185]=-38;
sine[9186]=-38;
sine[9187]=-38;
sine[9188]=-38;
sine[9189]=-38;
sine[9190]=-38;
sine[9191]=-38;
sine[9192]=-38;
sine[9193]=-38;
sine[9194]=-38;
sine[9195]=-38;
sine[9196]=-38;
sine[9197]=-38;
sine[9198]=-38;
sine[9199]=-38;
sine[9200]=-38;
sine[9201]=-38;
sine[9202]=-38;
sine[9203]=-38;
sine[9204]=-37;
sine[9205]=-37;
sine[9206]=-37;
sine[9207]=-37;
sine[9208]=-37;
sine[9209]=-37;
sine[9210]=-37;
sine[9211]=-37;
sine[9212]=-37;
sine[9213]=-37;
sine[9214]=-37;
sine[9215]=-37;
sine[9216]=-37;
sine[9217]=-37;
sine[9218]=-37;
sine[9219]=-37;
sine[9220]=-37;
sine[9221]=-37;
sine[9222]=-37;
sine[9223]=-37;
sine[9224]=-37;
sine[9225]=-37;
sine[9226]=-37;
sine[9227]=-36;
sine[9228]=-36;
sine[9229]=-36;
sine[9230]=-36;
sine[9231]=-36;
sine[9232]=-36;
sine[9233]=-36;
sine[9234]=-36;
sine[9235]=-36;
sine[9236]=-36;
sine[9237]=-36;
sine[9238]=-36;
sine[9239]=-36;
sine[9240]=-36;
sine[9241]=-36;
sine[9242]=-36;
sine[9243]=-36;
sine[9244]=-36;
sine[9245]=-36;
sine[9246]=-36;
sine[9247]=-36;
sine[9248]=-36;
sine[9249]=-36;
sine[9250]=-35;
sine[9251]=-35;
sine[9252]=-35;
sine[9253]=-35;
sine[9254]=-35;
sine[9255]=-35;
sine[9256]=-35;
sine[9257]=-35;
sine[9258]=-35;
sine[9259]=-35;
sine[9260]=-35;
sine[9261]=-35;
sine[9262]=-35;
sine[9263]=-35;
sine[9264]=-35;
sine[9265]=-35;
sine[9266]=-35;
sine[9267]=-35;
sine[9268]=-35;
sine[9269]=-35;
sine[9270]=-35;
sine[9271]=-35;
sine[9272]=-35;
sine[9273]=-34;
sine[9274]=-34;
sine[9275]=-34;
sine[9276]=-34;
sine[9277]=-34;
sine[9278]=-34;
sine[9279]=-34;
sine[9280]=-34;
sine[9281]=-34;
sine[9282]=-34;
sine[9283]=-34;
sine[9284]=-34;
sine[9285]=-34;
sine[9286]=-34;
sine[9287]=-34;
sine[9288]=-34;
sine[9289]=-34;
sine[9290]=-34;
sine[9291]=-34;
sine[9292]=-34;
sine[9293]=-34;
sine[9294]=-34;
sine[9295]=-33;
sine[9296]=-33;
sine[9297]=-33;
sine[9298]=-33;
sine[9299]=-33;
sine[9300]=-33;
sine[9301]=-33;
sine[9302]=-33;
sine[9303]=-33;
sine[9304]=-33;
sine[9305]=-33;
sine[9306]=-33;
sine[9307]=-33;
sine[9308]=-33;
sine[9309]=-33;
sine[9310]=-33;
sine[9311]=-33;
sine[9312]=-33;
sine[9313]=-33;
sine[9314]=-33;
sine[9315]=-33;
sine[9316]=-33;
sine[9317]=-33;
sine[9318]=-32;
sine[9319]=-32;
sine[9320]=-32;
sine[9321]=-32;
sine[9322]=-32;
sine[9323]=-32;
sine[9324]=-32;
sine[9325]=-32;
sine[9326]=-32;
sine[9327]=-32;
sine[9328]=-32;
sine[9329]=-32;
sine[9330]=-32;
sine[9331]=-32;
sine[9332]=-32;
sine[9333]=-32;
sine[9334]=-32;
sine[9335]=-32;
sine[9336]=-32;
sine[9337]=-32;
sine[9338]=-32;
sine[9339]=-32;
sine[9340]=-31;
sine[9341]=-31;
sine[9342]=-31;
sine[9343]=-31;
sine[9344]=-31;
sine[9345]=-31;
sine[9346]=-31;
sine[9347]=-31;
sine[9348]=-31;
sine[9349]=-31;
sine[9350]=-31;
sine[9351]=-31;
sine[9352]=-31;
sine[9353]=-31;
sine[9354]=-31;
sine[9355]=-31;
sine[9356]=-31;
sine[9357]=-31;
sine[9358]=-31;
sine[9359]=-31;
sine[9360]=-31;
sine[9361]=-31;
sine[9362]=-30;
sine[9363]=-30;
sine[9364]=-30;
sine[9365]=-30;
sine[9366]=-30;
sine[9367]=-30;
sine[9368]=-30;
sine[9369]=-30;
sine[9370]=-30;
sine[9371]=-30;
sine[9372]=-30;
sine[9373]=-30;
sine[9374]=-30;
sine[9375]=-30;
sine[9376]=-30;
sine[9377]=-30;
sine[9378]=-30;
sine[9379]=-30;
sine[9380]=-30;
sine[9381]=-30;
sine[9382]=-30;
sine[9383]=-30;
sine[9384]=-29;
sine[9385]=-29;
sine[9386]=-29;
sine[9387]=-29;
sine[9388]=-29;
sine[9389]=-29;
sine[9390]=-29;
sine[9391]=-29;
sine[9392]=-29;
sine[9393]=-29;
sine[9394]=-29;
sine[9395]=-29;
sine[9396]=-29;
sine[9397]=-29;
sine[9398]=-29;
sine[9399]=-29;
sine[9400]=-29;
sine[9401]=-29;
sine[9402]=-29;
sine[9403]=-29;
sine[9404]=-29;
sine[9405]=-29;
sine[9406]=-28;
sine[9407]=-28;
sine[9408]=-28;
sine[9409]=-28;
sine[9410]=-28;
sine[9411]=-28;
sine[9412]=-28;
sine[9413]=-28;
sine[9414]=-28;
sine[9415]=-28;
sine[9416]=-28;
sine[9417]=-28;
sine[9418]=-28;
sine[9419]=-28;
sine[9420]=-28;
sine[9421]=-28;
sine[9422]=-28;
sine[9423]=-28;
sine[9424]=-28;
sine[9425]=-28;
sine[9426]=-28;
sine[9427]=-28;
sine[9428]=-27;
sine[9429]=-27;
sine[9430]=-27;
sine[9431]=-27;
sine[9432]=-27;
sine[9433]=-27;
sine[9434]=-27;
sine[9435]=-27;
sine[9436]=-27;
sine[9437]=-27;
sine[9438]=-27;
sine[9439]=-27;
sine[9440]=-27;
sine[9441]=-27;
sine[9442]=-27;
sine[9443]=-27;
sine[9444]=-27;
sine[9445]=-27;
sine[9446]=-27;
sine[9447]=-27;
sine[9448]=-27;
sine[9449]=-27;
sine[9450]=-26;
sine[9451]=-26;
sine[9452]=-26;
sine[9453]=-26;
sine[9454]=-26;
sine[9455]=-26;
sine[9456]=-26;
sine[9457]=-26;
sine[9458]=-26;
sine[9459]=-26;
sine[9460]=-26;
sine[9461]=-26;
sine[9462]=-26;
sine[9463]=-26;
sine[9464]=-26;
sine[9465]=-26;
sine[9466]=-26;
sine[9467]=-26;
sine[9468]=-26;
sine[9469]=-26;
sine[9470]=-26;
sine[9471]=-25;
sine[9472]=-25;
sine[9473]=-25;
sine[9474]=-25;
sine[9475]=-25;
sine[9476]=-25;
sine[9477]=-25;
sine[9478]=-25;
sine[9479]=-25;
sine[9480]=-25;
sine[9481]=-25;
sine[9482]=-25;
sine[9483]=-25;
sine[9484]=-25;
sine[9485]=-25;
sine[9486]=-25;
sine[9487]=-25;
sine[9488]=-25;
sine[9489]=-25;
sine[9490]=-25;
sine[9491]=-25;
sine[9492]=-25;
sine[9493]=-24;
sine[9494]=-24;
sine[9495]=-24;
sine[9496]=-24;
sine[9497]=-24;
sine[9498]=-24;
sine[9499]=-24;
sine[9500]=-24;
sine[9501]=-24;
sine[9502]=-24;
sine[9503]=-24;
sine[9504]=-24;
sine[9505]=-24;
sine[9506]=-24;
sine[9507]=-24;
sine[9508]=-24;
sine[9509]=-24;
sine[9510]=-24;
sine[9511]=-24;
sine[9512]=-24;
sine[9513]=-24;
sine[9514]=-23;
sine[9515]=-23;
sine[9516]=-23;
sine[9517]=-23;
sine[9518]=-23;
sine[9519]=-23;
sine[9520]=-23;
sine[9521]=-23;
sine[9522]=-23;
sine[9523]=-23;
sine[9524]=-23;
sine[9525]=-23;
sine[9526]=-23;
sine[9527]=-23;
sine[9528]=-23;
sine[9529]=-23;
sine[9530]=-23;
sine[9531]=-23;
sine[9532]=-23;
sine[9533]=-23;
sine[9534]=-23;
sine[9535]=-23;
sine[9536]=-22;
sine[9537]=-22;
sine[9538]=-22;
sine[9539]=-22;
sine[9540]=-22;
sine[9541]=-22;
sine[9542]=-22;
sine[9543]=-22;
sine[9544]=-22;
sine[9545]=-22;
sine[9546]=-22;
sine[9547]=-22;
sine[9548]=-22;
sine[9549]=-22;
sine[9550]=-22;
sine[9551]=-22;
sine[9552]=-22;
sine[9553]=-22;
sine[9554]=-22;
sine[9555]=-22;
sine[9556]=-22;
sine[9557]=-21;
sine[9558]=-21;
sine[9559]=-21;
sine[9560]=-21;
sine[9561]=-21;
sine[9562]=-21;
sine[9563]=-21;
sine[9564]=-21;
sine[9565]=-21;
sine[9566]=-21;
sine[9567]=-21;
sine[9568]=-21;
sine[9569]=-21;
sine[9570]=-21;
sine[9571]=-21;
sine[9572]=-21;
sine[9573]=-21;
sine[9574]=-21;
sine[9575]=-21;
sine[9576]=-21;
sine[9577]=-21;
sine[9578]=-20;
sine[9579]=-20;
sine[9580]=-20;
sine[9581]=-20;
sine[9582]=-20;
sine[9583]=-20;
sine[9584]=-20;
sine[9585]=-20;
sine[9586]=-20;
sine[9587]=-20;
sine[9588]=-20;
sine[9589]=-20;
sine[9590]=-20;
sine[9591]=-20;
sine[9592]=-20;
sine[9593]=-20;
sine[9594]=-20;
sine[9595]=-20;
sine[9596]=-20;
sine[9597]=-20;
sine[9598]=-20;
sine[9599]=-19;
sine[9600]=-19;
sine[9601]=-19;
sine[9602]=-19;
sine[9603]=-19;
sine[9604]=-19;
sine[9605]=-19;
sine[9606]=-19;
sine[9607]=-19;
sine[9608]=-19;
sine[9609]=-19;
sine[9610]=-19;
sine[9611]=-19;
sine[9612]=-19;
sine[9613]=-19;
sine[9614]=-19;
sine[9615]=-19;
sine[9616]=-19;
sine[9617]=-19;
sine[9618]=-19;
sine[9619]=-19;
sine[9620]=-18;
sine[9621]=-18;
sine[9622]=-18;
sine[9623]=-18;
sine[9624]=-18;
sine[9625]=-18;
sine[9626]=-18;
sine[9627]=-18;
sine[9628]=-18;
sine[9629]=-18;
sine[9630]=-18;
sine[9631]=-18;
sine[9632]=-18;
sine[9633]=-18;
sine[9634]=-18;
sine[9635]=-18;
sine[9636]=-18;
sine[9637]=-18;
sine[9638]=-18;
sine[9639]=-18;
sine[9640]=-18;
sine[9641]=-17;
sine[9642]=-17;
sine[9643]=-17;
sine[9644]=-17;
sine[9645]=-17;
sine[9646]=-17;
sine[9647]=-17;
sine[9648]=-17;
sine[9649]=-17;
sine[9650]=-17;
sine[9651]=-17;
sine[9652]=-17;
sine[9653]=-17;
sine[9654]=-17;
sine[9655]=-17;
sine[9656]=-17;
sine[9657]=-17;
sine[9658]=-17;
sine[9659]=-17;
sine[9660]=-17;
sine[9661]=-17;
sine[9662]=-16;
sine[9663]=-16;
sine[9664]=-16;
sine[9665]=-16;
sine[9666]=-16;
sine[9667]=-16;
sine[9668]=-16;
sine[9669]=-16;
sine[9670]=-16;
sine[9671]=-16;
sine[9672]=-16;
sine[9673]=-16;
sine[9674]=-16;
sine[9675]=-16;
sine[9676]=-16;
sine[9677]=-16;
sine[9678]=-16;
sine[9679]=-16;
sine[9680]=-16;
sine[9681]=-16;
sine[9682]=-16;
sine[9683]=-15;
sine[9684]=-15;
sine[9685]=-15;
sine[9686]=-15;
sine[9687]=-15;
sine[9688]=-15;
sine[9689]=-15;
sine[9690]=-15;
sine[9691]=-15;
sine[9692]=-15;
sine[9693]=-15;
sine[9694]=-15;
sine[9695]=-15;
sine[9696]=-15;
sine[9697]=-15;
sine[9698]=-15;
sine[9699]=-15;
sine[9700]=-15;
sine[9701]=-15;
sine[9702]=-15;
sine[9703]=-14;
sine[9704]=-14;
sine[9705]=-14;
sine[9706]=-14;
sine[9707]=-14;
sine[9708]=-14;
sine[9709]=-14;
sine[9710]=-14;
sine[9711]=-14;
sine[9712]=-14;
sine[9713]=-14;
sine[9714]=-14;
sine[9715]=-14;
sine[9716]=-14;
sine[9717]=-14;
sine[9718]=-14;
sine[9719]=-14;
sine[9720]=-14;
sine[9721]=-14;
sine[9722]=-14;
sine[9723]=-14;
sine[9724]=-13;
sine[9725]=-13;
sine[9726]=-13;
sine[9727]=-13;
sine[9728]=-13;
sine[9729]=-13;
sine[9730]=-13;
sine[9731]=-13;
sine[9732]=-13;
sine[9733]=-13;
sine[9734]=-13;
sine[9735]=-13;
sine[9736]=-13;
sine[9737]=-13;
sine[9738]=-13;
sine[9739]=-13;
sine[9740]=-13;
sine[9741]=-13;
sine[9742]=-13;
sine[9743]=-13;
sine[9744]=-13;
sine[9745]=-12;
sine[9746]=-12;
sine[9747]=-12;
sine[9748]=-12;
sine[9749]=-12;
sine[9750]=-12;
sine[9751]=-12;
sine[9752]=-12;
sine[9753]=-12;
sine[9754]=-12;
sine[9755]=-12;
sine[9756]=-12;
sine[9757]=-12;
sine[9758]=-12;
sine[9759]=-12;
sine[9760]=-12;
sine[9761]=-12;
sine[9762]=-12;
sine[9763]=-12;
sine[9764]=-12;
sine[9765]=-11;
sine[9766]=-11;
sine[9767]=-11;
sine[9768]=-11;
sine[9769]=-11;
sine[9770]=-11;
sine[9771]=-11;
sine[9772]=-11;
sine[9773]=-11;
sine[9774]=-11;
sine[9775]=-11;
sine[9776]=-11;
sine[9777]=-11;
sine[9778]=-11;
sine[9779]=-11;
sine[9780]=-11;
sine[9781]=-11;
sine[9782]=-11;
sine[9783]=-11;
sine[9784]=-11;
sine[9785]=-11;
sine[9786]=-10;
sine[9787]=-10;
sine[9788]=-10;
sine[9789]=-10;
sine[9790]=-10;
sine[9791]=-10;
sine[9792]=-10;
sine[9793]=-10;
sine[9794]=-10;
sine[9795]=-10;
sine[9796]=-10;
sine[9797]=-10;
sine[9798]=-10;
sine[9799]=-10;
sine[9800]=-10;
sine[9801]=-10;
sine[9802]=-10;
sine[9803]=-10;
sine[9804]=-10;
sine[9805]=-10;
sine[9806]=-9;
sine[9807]=-9;
sine[9808]=-9;
sine[9809]=-9;
sine[9810]=-9;
sine[9811]=-9;
sine[9812]=-9;
sine[9813]=-9;
sine[9814]=-9;
sine[9815]=-9;
sine[9816]=-9;
sine[9817]=-9;
sine[9818]=-9;
sine[9819]=-9;
sine[9820]=-9;
sine[9821]=-9;
sine[9822]=-9;
sine[9823]=-9;
sine[9824]=-9;
sine[9825]=-9;
sine[9826]=-9;
sine[9827]=-8;
sine[9828]=-8;
sine[9829]=-8;
sine[9830]=-8;
sine[9831]=-8;
sine[9832]=-8;
sine[9833]=-8;
sine[9834]=-8;
sine[9835]=-8;
sine[9836]=-8;
sine[9837]=-8;
sine[9838]=-8;
sine[9839]=-8;
sine[9840]=-8;
sine[9841]=-8;
sine[9842]=-8;
sine[9843]=-8;
sine[9844]=-8;
sine[9845]=-8;
sine[9846]=-8;
sine[9847]=-7;
sine[9848]=-7;
sine[9849]=-7;
sine[9850]=-7;
sine[9851]=-7;
sine[9852]=-7;
sine[9853]=-7;
sine[9854]=-7;
sine[9855]=-7;
sine[9856]=-7;
sine[9857]=-7;
sine[9858]=-7;
sine[9859]=-7;
sine[9860]=-7;
sine[9861]=-7;
sine[9862]=-7;
sine[9863]=-7;
sine[9864]=-7;
sine[9865]=-7;
sine[9866]=-7;
sine[9867]=-7;
sine[9868]=-6;
sine[9869]=-6;
sine[9870]=-6;
sine[9871]=-6;
sine[9872]=-6;
sine[9873]=-6;
sine[9874]=-6;
sine[9875]=-6;
sine[9876]=-6;
sine[9877]=-6;
sine[9878]=-6;
sine[9879]=-6;
sine[9880]=-6;
sine[9881]=-6;
sine[9882]=-6;
sine[9883]=-6;
sine[9884]=-6;
sine[9885]=-6;
sine[9886]=-6;
sine[9887]=-6;
sine[9888]=-5;
sine[9889]=-5;
sine[9890]=-5;
sine[9891]=-5;
sine[9892]=-5;
sine[9893]=-5;
sine[9894]=-5;
sine[9895]=-5;
sine[9896]=-5;
sine[9897]=-5;
sine[9898]=-5;
sine[9899]=-5;
sine[9900]=-5;
sine[9901]=-5;
sine[9902]=-5;
sine[9903]=-5;
sine[9904]=-5;
sine[9905]=-5;
sine[9906]=-5;
sine[9907]=-5;
sine[9908]=-5;
sine[9909]=-4;
sine[9910]=-4;
sine[9911]=-4;
sine[9912]=-4;
sine[9913]=-4;
sine[9914]=-4;
sine[9915]=-4;
sine[9916]=-4;
sine[9917]=-4;
sine[9918]=-4;
sine[9919]=-4;
sine[9920]=-4;
sine[9921]=-4;
sine[9922]=-4;
sine[9923]=-4;
sine[9924]=-4;
sine[9925]=-4;
sine[9926]=-4;
sine[9927]=-4;
sine[9928]=-4;
sine[9929]=-3;
sine[9930]=-3;
sine[9931]=-3;
sine[9932]=-3;
sine[9933]=-3;
sine[9934]=-3;
sine[9935]=-3;
sine[9936]=-3;
sine[9937]=-3;
sine[9938]=-3;
sine[9939]=-3;
sine[9940]=-3;
sine[9941]=-3;
sine[9942]=-3;
sine[9943]=-3;
sine[9944]=-3;
sine[9945]=-3;
sine[9946]=-3;
sine[9947]=-3;
sine[9948]=-3;
sine[9949]=-3;
sine[9950]=-2;
sine[9951]=-2;
sine[9952]=-2;
sine[9953]=-2;
sine[9954]=-2;
sine[9955]=-2;
sine[9956]=-2;
sine[9957]=-2;
sine[9958]=-2;
sine[9959]=-2;
sine[9960]=-2;
sine[9961]=-2;
sine[9962]=-2;
sine[9963]=-2;
sine[9964]=-2;
sine[9965]=-2;
sine[9966]=-2;
sine[9967]=-2;
sine[9968]=-2;
sine[9969]=-2;
sine[9970]=-1;
sine[9971]=-1;
sine[9972]=-1;
sine[9973]=-1;
sine[9974]=-1;
sine[9975]=-1;
sine[9976]=-1;
sine[9977]=-1;
sine[9978]=-1;
sine[9979]=-1;
sine[9980]=-1;
sine[9981]=-1;
sine[9982]=-1;
sine[9983]=-1;
sine[9984]=-1;
sine[9985]=-1;
sine[9986]=-1;
sine[9987]=-1;
sine[9988]=-1;
sine[9989]=-1;
sine[9990]=0;
sine[9991]=0;
sine[9992]=0;
sine[9993]=0;
sine[9994]=0;
sine[9995]=0;
sine[9996]=0;
sine[9997]=0;
sine[9998]=0;
sine[9999]=0;
sine[10000]=0;
sine[10001]=0;
sine[10002]=0;
sine[10003]=0;
sine[10004]=0;
sine[10005]=0;
sine[10006]=0;
sine[10007]=0;
sine[10008]=0;
sine[10009]=0;
sine[10010]=0;
sine[10011]=1;
sine[10012]=1;
sine[10013]=1;
sine[10014]=1;
sine[10015]=1;
sine[10016]=1;
sine[10017]=1;
sine[10018]=1;
sine[10019]=1;
sine[10020]=1;
sine[10021]=1;
sine[10022]=1;
sine[10023]=1;
sine[10024]=1;
sine[10025]=1;
sine[10026]=1;
sine[10027]=1;
sine[10028]=1;
sine[10029]=1;
sine[10030]=1;
sine[10031]=2;
sine[10032]=2;
sine[10033]=2;
sine[10034]=2;
sine[10035]=2;
sine[10036]=2;
sine[10037]=2;
sine[10038]=2;
sine[10039]=2;
sine[10040]=2;
sine[10041]=2;
sine[10042]=2;
sine[10043]=2;
sine[10044]=2;
sine[10045]=2;
sine[10046]=2;
sine[10047]=2;
sine[10048]=2;
sine[10049]=2;
sine[10050]=2;
sine[10051]=3;
sine[10052]=3;
sine[10053]=3;
sine[10054]=3;
sine[10055]=3;
sine[10056]=3;
sine[10057]=3;
sine[10058]=3;
sine[10059]=3;
sine[10060]=3;
sine[10061]=3;
sine[10062]=3;
sine[10063]=3;
sine[10064]=3;
sine[10065]=3;
sine[10066]=3;
sine[10067]=3;
sine[10068]=3;
sine[10069]=3;
sine[10070]=3;
sine[10071]=3;
sine[10072]=4;
sine[10073]=4;
sine[10074]=4;
sine[10075]=4;
sine[10076]=4;
sine[10077]=4;
sine[10078]=4;
sine[10079]=4;
sine[10080]=4;
sine[10081]=4;
sine[10082]=4;
sine[10083]=4;
sine[10084]=4;
sine[10085]=4;
sine[10086]=4;
sine[10087]=4;
sine[10088]=4;
sine[10089]=4;
sine[10090]=4;
sine[10091]=4;
sine[10092]=5;
sine[10093]=5;
sine[10094]=5;
sine[10095]=5;
sine[10096]=5;
sine[10097]=5;
sine[10098]=5;
sine[10099]=5;
sine[10100]=5;
sine[10101]=5;
sine[10102]=5;
sine[10103]=5;
sine[10104]=5;
sine[10105]=5;
sine[10106]=5;
sine[10107]=5;
sine[10108]=5;
sine[10109]=5;
sine[10110]=5;
sine[10111]=5;
sine[10112]=5;
sine[10113]=6;
sine[10114]=6;
sine[10115]=6;
sine[10116]=6;
sine[10117]=6;
sine[10118]=6;
sine[10119]=6;
sine[10120]=6;
sine[10121]=6;
sine[10122]=6;
sine[10123]=6;
sine[10124]=6;
sine[10125]=6;
sine[10126]=6;
sine[10127]=6;
sine[10128]=6;
sine[10129]=6;
sine[10130]=6;
sine[10131]=6;
sine[10132]=6;
sine[10133]=7;
sine[10134]=7;
sine[10135]=7;
sine[10136]=7;
sine[10137]=7;
sine[10138]=7;
sine[10139]=7;
sine[10140]=7;
sine[10141]=7;
sine[10142]=7;
sine[10143]=7;
sine[10144]=7;
sine[10145]=7;
sine[10146]=7;
sine[10147]=7;
sine[10148]=7;
sine[10149]=7;
sine[10150]=7;
sine[10151]=7;
sine[10152]=7;
sine[10153]=7;
sine[10154]=8;
sine[10155]=8;
sine[10156]=8;
sine[10157]=8;
sine[10158]=8;
sine[10159]=8;
sine[10160]=8;
sine[10161]=8;
sine[10162]=8;
sine[10163]=8;
sine[10164]=8;
sine[10165]=8;
sine[10166]=8;
sine[10167]=8;
sine[10168]=8;
sine[10169]=8;
sine[10170]=8;
sine[10171]=8;
sine[10172]=8;
sine[10173]=8;
sine[10174]=9;
sine[10175]=9;
sine[10176]=9;
sine[10177]=9;
sine[10178]=9;
sine[10179]=9;
sine[10180]=9;
sine[10181]=9;
sine[10182]=9;
sine[10183]=9;
sine[10184]=9;
sine[10185]=9;
sine[10186]=9;
sine[10187]=9;
sine[10188]=9;
sine[10189]=9;
sine[10190]=9;
sine[10191]=9;
sine[10192]=9;
sine[10193]=9;
sine[10194]=9;
sine[10195]=10;
sine[10196]=10;
sine[10197]=10;
sine[10198]=10;
sine[10199]=10;
sine[10200]=10;
sine[10201]=10;
sine[10202]=10;
sine[10203]=10;
sine[10204]=10;
sine[10205]=10;
sine[10206]=10;
sine[10207]=10;
sine[10208]=10;
sine[10209]=10;
sine[10210]=10;
sine[10211]=10;
sine[10212]=10;
sine[10213]=10;
sine[10214]=10;
sine[10215]=11;
sine[10216]=11;
sine[10217]=11;
sine[10218]=11;
sine[10219]=11;
sine[10220]=11;
sine[10221]=11;
sine[10222]=11;
sine[10223]=11;
sine[10224]=11;
sine[10225]=11;
sine[10226]=11;
sine[10227]=11;
sine[10228]=11;
sine[10229]=11;
sine[10230]=11;
sine[10231]=11;
sine[10232]=11;
sine[10233]=11;
sine[10234]=11;
sine[10235]=11;
sine[10236]=12;
sine[10237]=12;
sine[10238]=12;
sine[10239]=12;
sine[10240]=12;
sine[10241]=12;
sine[10242]=12;
sine[10243]=12;
sine[10244]=12;
sine[10245]=12;
sine[10246]=12;
sine[10247]=12;
sine[10248]=12;
sine[10249]=12;
sine[10250]=12;
sine[10251]=12;
sine[10252]=12;
sine[10253]=12;
sine[10254]=12;
sine[10255]=12;
sine[10256]=13;
sine[10257]=13;
sine[10258]=13;
sine[10259]=13;
sine[10260]=13;
sine[10261]=13;
sine[10262]=13;
sine[10263]=13;
sine[10264]=13;
sine[10265]=13;
sine[10266]=13;
sine[10267]=13;
sine[10268]=13;
sine[10269]=13;
sine[10270]=13;
sine[10271]=13;
sine[10272]=13;
sine[10273]=13;
sine[10274]=13;
sine[10275]=13;
sine[10276]=13;
sine[10277]=14;
sine[10278]=14;
sine[10279]=14;
sine[10280]=14;
sine[10281]=14;
sine[10282]=14;
sine[10283]=14;
sine[10284]=14;
sine[10285]=14;
sine[10286]=14;
sine[10287]=14;
sine[10288]=14;
sine[10289]=14;
sine[10290]=14;
sine[10291]=14;
sine[10292]=14;
sine[10293]=14;
sine[10294]=14;
sine[10295]=14;
sine[10296]=14;
sine[10297]=14;
sine[10298]=15;
sine[10299]=15;
sine[10300]=15;
sine[10301]=15;
sine[10302]=15;
sine[10303]=15;
sine[10304]=15;
sine[10305]=15;
sine[10306]=15;
sine[10307]=15;
sine[10308]=15;
sine[10309]=15;
sine[10310]=15;
sine[10311]=15;
sine[10312]=15;
sine[10313]=15;
sine[10314]=15;
sine[10315]=15;
sine[10316]=15;
sine[10317]=15;
sine[10318]=16;
sine[10319]=16;
sine[10320]=16;
sine[10321]=16;
sine[10322]=16;
sine[10323]=16;
sine[10324]=16;
sine[10325]=16;
sine[10326]=16;
sine[10327]=16;
sine[10328]=16;
sine[10329]=16;
sine[10330]=16;
sine[10331]=16;
sine[10332]=16;
sine[10333]=16;
sine[10334]=16;
sine[10335]=16;
sine[10336]=16;
sine[10337]=16;
sine[10338]=16;
sine[10339]=17;
sine[10340]=17;
sine[10341]=17;
sine[10342]=17;
sine[10343]=17;
sine[10344]=17;
sine[10345]=17;
sine[10346]=17;
sine[10347]=17;
sine[10348]=17;
sine[10349]=17;
sine[10350]=17;
sine[10351]=17;
sine[10352]=17;
sine[10353]=17;
sine[10354]=17;
sine[10355]=17;
sine[10356]=17;
sine[10357]=17;
sine[10358]=17;
sine[10359]=17;
sine[10360]=18;
sine[10361]=18;
sine[10362]=18;
sine[10363]=18;
sine[10364]=18;
sine[10365]=18;
sine[10366]=18;
sine[10367]=18;
sine[10368]=18;
sine[10369]=18;
sine[10370]=18;
sine[10371]=18;
sine[10372]=18;
sine[10373]=18;
sine[10374]=18;
sine[10375]=18;
sine[10376]=18;
sine[10377]=18;
sine[10378]=18;
sine[10379]=18;
sine[10380]=18;
sine[10381]=19;
sine[10382]=19;
sine[10383]=19;
sine[10384]=19;
sine[10385]=19;
sine[10386]=19;
sine[10387]=19;
sine[10388]=19;
sine[10389]=19;
sine[10390]=19;
sine[10391]=19;
sine[10392]=19;
sine[10393]=19;
sine[10394]=19;
sine[10395]=19;
sine[10396]=19;
sine[10397]=19;
sine[10398]=19;
sine[10399]=19;
sine[10400]=19;
sine[10401]=19;
sine[10402]=20;
sine[10403]=20;
sine[10404]=20;
sine[10405]=20;
sine[10406]=20;
sine[10407]=20;
sine[10408]=20;
sine[10409]=20;
sine[10410]=20;
sine[10411]=20;
sine[10412]=20;
sine[10413]=20;
sine[10414]=20;
sine[10415]=20;
sine[10416]=20;
sine[10417]=20;
sine[10418]=20;
sine[10419]=20;
sine[10420]=20;
sine[10421]=20;
sine[10422]=20;
sine[10423]=21;
sine[10424]=21;
sine[10425]=21;
sine[10426]=21;
sine[10427]=21;
sine[10428]=21;
sine[10429]=21;
sine[10430]=21;
sine[10431]=21;
sine[10432]=21;
sine[10433]=21;
sine[10434]=21;
sine[10435]=21;
sine[10436]=21;
sine[10437]=21;
sine[10438]=21;
sine[10439]=21;
sine[10440]=21;
sine[10441]=21;
sine[10442]=21;
sine[10443]=21;
sine[10444]=22;
sine[10445]=22;
sine[10446]=22;
sine[10447]=22;
sine[10448]=22;
sine[10449]=22;
sine[10450]=22;
sine[10451]=22;
sine[10452]=22;
sine[10453]=22;
sine[10454]=22;
sine[10455]=22;
sine[10456]=22;
sine[10457]=22;
sine[10458]=22;
sine[10459]=22;
sine[10460]=22;
sine[10461]=22;
sine[10462]=22;
sine[10463]=22;
sine[10464]=22;
sine[10465]=23;
sine[10466]=23;
sine[10467]=23;
sine[10468]=23;
sine[10469]=23;
sine[10470]=23;
sine[10471]=23;
sine[10472]=23;
sine[10473]=23;
sine[10474]=23;
sine[10475]=23;
sine[10476]=23;
sine[10477]=23;
sine[10478]=23;
sine[10479]=23;
sine[10480]=23;
sine[10481]=23;
sine[10482]=23;
sine[10483]=23;
sine[10484]=23;
sine[10485]=23;
sine[10486]=23;
sine[10487]=24;
sine[10488]=24;
sine[10489]=24;
sine[10490]=24;
sine[10491]=24;
sine[10492]=24;
sine[10493]=24;
sine[10494]=24;
sine[10495]=24;
sine[10496]=24;
sine[10497]=24;
sine[10498]=24;
sine[10499]=24;
sine[10500]=24;
sine[10501]=24;
sine[10502]=24;
sine[10503]=24;
sine[10504]=24;
sine[10505]=24;
sine[10506]=24;
sine[10507]=24;
sine[10508]=25;
sine[10509]=25;
sine[10510]=25;
sine[10511]=25;
sine[10512]=25;
sine[10513]=25;
sine[10514]=25;
sine[10515]=25;
sine[10516]=25;
sine[10517]=25;
sine[10518]=25;
sine[10519]=25;
sine[10520]=25;
sine[10521]=25;
sine[10522]=25;
sine[10523]=25;
sine[10524]=25;
sine[10525]=25;
sine[10526]=25;
sine[10527]=25;
sine[10528]=25;
sine[10529]=25;
sine[10530]=26;
sine[10531]=26;
sine[10532]=26;
sine[10533]=26;
sine[10534]=26;
sine[10535]=26;
sine[10536]=26;
sine[10537]=26;
sine[10538]=26;
sine[10539]=26;
sine[10540]=26;
sine[10541]=26;
sine[10542]=26;
sine[10543]=26;
sine[10544]=26;
sine[10545]=26;
sine[10546]=26;
sine[10547]=26;
sine[10548]=26;
sine[10549]=26;
sine[10550]=26;
sine[10551]=27;
sine[10552]=27;
sine[10553]=27;
sine[10554]=27;
sine[10555]=27;
sine[10556]=27;
sine[10557]=27;
sine[10558]=27;
sine[10559]=27;
sine[10560]=27;
sine[10561]=27;
sine[10562]=27;
sine[10563]=27;
sine[10564]=27;
sine[10565]=27;
sine[10566]=27;
sine[10567]=27;
sine[10568]=27;
sine[10569]=27;
sine[10570]=27;
sine[10571]=27;
sine[10572]=27;
sine[10573]=28;
sine[10574]=28;
sine[10575]=28;
sine[10576]=28;
sine[10577]=28;
sine[10578]=28;
sine[10579]=28;
sine[10580]=28;
sine[10581]=28;
sine[10582]=28;
sine[10583]=28;
sine[10584]=28;
sine[10585]=28;
sine[10586]=28;
sine[10587]=28;
sine[10588]=28;
sine[10589]=28;
sine[10590]=28;
sine[10591]=28;
sine[10592]=28;
sine[10593]=28;
sine[10594]=28;
sine[10595]=29;
sine[10596]=29;
sine[10597]=29;
sine[10598]=29;
sine[10599]=29;
sine[10600]=29;
sine[10601]=29;
sine[10602]=29;
sine[10603]=29;
sine[10604]=29;
sine[10605]=29;
sine[10606]=29;
sine[10607]=29;
sine[10608]=29;
sine[10609]=29;
sine[10610]=29;
sine[10611]=29;
sine[10612]=29;
sine[10613]=29;
sine[10614]=29;
sine[10615]=29;
sine[10616]=29;
sine[10617]=30;
sine[10618]=30;
sine[10619]=30;
sine[10620]=30;
sine[10621]=30;
sine[10622]=30;
sine[10623]=30;
sine[10624]=30;
sine[10625]=30;
sine[10626]=30;
sine[10627]=30;
sine[10628]=30;
sine[10629]=30;
sine[10630]=30;
sine[10631]=30;
sine[10632]=30;
sine[10633]=30;
sine[10634]=30;
sine[10635]=30;
sine[10636]=30;
sine[10637]=30;
sine[10638]=30;
sine[10639]=31;
sine[10640]=31;
sine[10641]=31;
sine[10642]=31;
sine[10643]=31;
sine[10644]=31;
sine[10645]=31;
sine[10646]=31;
sine[10647]=31;
sine[10648]=31;
sine[10649]=31;
sine[10650]=31;
sine[10651]=31;
sine[10652]=31;
sine[10653]=31;
sine[10654]=31;
sine[10655]=31;
sine[10656]=31;
sine[10657]=31;
sine[10658]=31;
sine[10659]=31;
sine[10660]=31;
sine[10661]=32;
sine[10662]=32;
sine[10663]=32;
sine[10664]=32;
sine[10665]=32;
sine[10666]=32;
sine[10667]=32;
sine[10668]=32;
sine[10669]=32;
sine[10670]=32;
sine[10671]=32;
sine[10672]=32;
sine[10673]=32;
sine[10674]=32;
sine[10675]=32;
sine[10676]=32;
sine[10677]=32;
sine[10678]=32;
sine[10679]=32;
sine[10680]=32;
sine[10681]=32;
sine[10682]=32;
sine[10683]=33;
sine[10684]=33;
sine[10685]=33;
sine[10686]=33;
sine[10687]=33;
sine[10688]=33;
sine[10689]=33;
sine[10690]=33;
sine[10691]=33;
sine[10692]=33;
sine[10693]=33;
sine[10694]=33;
sine[10695]=33;
sine[10696]=33;
sine[10697]=33;
sine[10698]=33;
sine[10699]=33;
sine[10700]=33;
sine[10701]=33;
sine[10702]=33;
sine[10703]=33;
sine[10704]=33;
sine[10705]=33;
sine[10706]=34;
sine[10707]=34;
sine[10708]=34;
sine[10709]=34;
sine[10710]=34;
sine[10711]=34;
sine[10712]=34;
sine[10713]=34;
sine[10714]=34;
sine[10715]=34;
sine[10716]=34;
sine[10717]=34;
sine[10718]=34;
sine[10719]=34;
sine[10720]=34;
sine[10721]=34;
sine[10722]=34;
sine[10723]=34;
sine[10724]=34;
sine[10725]=34;
sine[10726]=34;
sine[10727]=34;
sine[10728]=35;
sine[10729]=35;
sine[10730]=35;
sine[10731]=35;
sine[10732]=35;
sine[10733]=35;
sine[10734]=35;
sine[10735]=35;
sine[10736]=35;
sine[10737]=35;
sine[10738]=35;
sine[10739]=35;
sine[10740]=35;
sine[10741]=35;
sine[10742]=35;
sine[10743]=35;
sine[10744]=35;
sine[10745]=35;
sine[10746]=35;
sine[10747]=35;
sine[10748]=35;
sine[10749]=35;
sine[10750]=35;
sine[10751]=36;
sine[10752]=36;
sine[10753]=36;
sine[10754]=36;
sine[10755]=36;
sine[10756]=36;
sine[10757]=36;
sine[10758]=36;
sine[10759]=36;
sine[10760]=36;
sine[10761]=36;
sine[10762]=36;
sine[10763]=36;
sine[10764]=36;
sine[10765]=36;
sine[10766]=36;
sine[10767]=36;
sine[10768]=36;
sine[10769]=36;
sine[10770]=36;
sine[10771]=36;
sine[10772]=36;
sine[10773]=36;
sine[10774]=37;
sine[10775]=37;
sine[10776]=37;
sine[10777]=37;
sine[10778]=37;
sine[10779]=37;
sine[10780]=37;
sine[10781]=37;
sine[10782]=37;
sine[10783]=37;
sine[10784]=37;
sine[10785]=37;
sine[10786]=37;
sine[10787]=37;
sine[10788]=37;
sine[10789]=37;
sine[10790]=37;
sine[10791]=37;
sine[10792]=37;
sine[10793]=37;
sine[10794]=37;
sine[10795]=37;
sine[10796]=37;
sine[10797]=38;
sine[10798]=38;
sine[10799]=38;
sine[10800]=38;
sine[10801]=38;
sine[10802]=38;
sine[10803]=38;
sine[10804]=38;
sine[10805]=38;
sine[10806]=38;
sine[10807]=38;
sine[10808]=38;
sine[10809]=38;
sine[10810]=38;
sine[10811]=38;
sine[10812]=38;
sine[10813]=38;
sine[10814]=38;
sine[10815]=38;
sine[10816]=38;
sine[10817]=38;
sine[10818]=38;
sine[10819]=38;
sine[10820]=38;
sine[10821]=39;
sine[10822]=39;
sine[10823]=39;
sine[10824]=39;
sine[10825]=39;
sine[10826]=39;
sine[10827]=39;
sine[10828]=39;
sine[10829]=39;
sine[10830]=39;
sine[10831]=39;
sine[10832]=39;
sine[10833]=39;
sine[10834]=39;
sine[10835]=39;
sine[10836]=39;
sine[10837]=39;
sine[10838]=39;
sine[10839]=39;
sine[10840]=39;
sine[10841]=39;
sine[10842]=39;
sine[10843]=39;
sine[10844]=40;
sine[10845]=40;
sine[10846]=40;
sine[10847]=40;
sine[10848]=40;
sine[10849]=40;
sine[10850]=40;
sine[10851]=40;
sine[10852]=40;
sine[10853]=40;
sine[10854]=40;
sine[10855]=40;
sine[10856]=40;
sine[10857]=40;
sine[10858]=40;
sine[10859]=40;
sine[10860]=40;
sine[10861]=40;
sine[10862]=40;
sine[10863]=40;
sine[10864]=40;
sine[10865]=40;
sine[10866]=40;
sine[10867]=40;
sine[10868]=41;
sine[10869]=41;
sine[10870]=41;
sine[10871]=41;
sine[10872]=41;
sine[10873]=41;
sine[10874]=41;
sine[10875]=41;
sine[10876]=41;
sine[10877]=41;
sine[10878]=41;
sine[10879]=41;
sine[10880]=41;
sine[10881]=41;
sine[10882]=41;
sine[10883]=41;
sine[10884]=41;
sine[10885]=41;
sine[10886]=41;
sine[10887]=41;
sine[10888]=41;
sine[10889]=41;
sine[10890]=41;
sine[10891]=41;
sine[10892]=42;
sine[10893]=42;
sine[10894]=42;
sine[10895]=42;
sine[10896]=42;
sine[10897]=42;
sine[10898]=42;
sine[10899]=42;
sine[10900]=42;
sine[10901]=42;
sine[10902]=42;
sine[10903]=42;
sine[10904]=42;
sine[10905]=42;
sine[10906]=42;
sine[10907]=42;
sine[10908]=42;
sine[10909]=42;
sine[10910]=42;
sine[10911]=42;
sine[10912]=42;
sine[10913]=42;
sine[10914]=42;
sine[10915]=42;
sine[10916]=43;
sine[10917]=43;
sine[10918]=43;
sine[10919]=43;
sine[10920]=43;
sine[10921]=43;
sine[10922]=43;
sine[10923]=43;
sine[10924]=43;
sine[10925]=43;
sine[10926]=43;
sine[10927]=43;
sine[10928]=43;
sine[10929]=43;
sine[10930]=43;
sine[10931]=43;
sine[10932]=43;
sine[10933]=43;
sine[10934]=43;
sine[10935]=43;
sine[10936]=43;
sine[10937]=43;
sine[10938]=43;
sine[10939]=43;
sine[10940]=44;
sine[10941]=44;
sine[10942]=44;
sine[10943]=44;
sine[10944]=44;
sine[10945]=44;
sine[10946]=44;
sine[10947]=44;
sine[10948]=44;
sine[10949]=44;
sine[10950]=44;
sine[10951]=44;
sine[10952]=44;
sine[10953]=44;
sine[10954]=44;
sine[10955]=44;
sine[10956]=44;
sine[10957]=44;
sine[10958]=44;
sine[10959]=44;
sine[10960]=44;
sine[10961]=44;
sine[10962]=44;
sine[10963]=44;
sine[10964]=44;
sine[10965]=45;
sine[10966]=45;
sine[10967]=45;
sine[10968]=45;
sine[10969]=45;
sine[10970]=45;
sine[10971]=45;
sine[10972]=45;
sine[10973]=45;
sine[10974]=45;
sine[10975]=45;
sine[10976]=45;
sine[10977]=45;
sine[10978]=45;
sine[10979]=45;
sine[10980]=45;
sine[10981]=45;
sine[10982]=45;
sine[10983]=45;
sine[10984]=45;
sine[10985]=45;
sine[10986]=45;
sine[10987]=45;
sine[10988]=45;
sine[10989]=45;
sine[10990]=46;
sine[10991]=46;
sine[10992]=46;
sine[10993]=46;
sine[10994]=46;
sine[10995]=46;
sine[10996]=46;
sine[10997]=46;
sine[10998]=46;
sine[10999]=46;
sine[11000]=46;
sine[11001]=46;
sine[11002]=46;
sine[11003]=46;
sine[11004]=46;
sine[11005]=46;
sine[11006]=46;
sine[11007]=46;
sine[11008]=46;
sine[11009]=46;
sine[11010]=46;
sine[11011]=46;
sine[11012]=46;
sine[11013]=46;
sine[11014]=46;
sine[11015]=47;
sine[11016]=47;
sine[11017]=47;
sine[11018]=47;
sine[11019]=47;
sine[11020]=47;
sine[11021]=47;
sine[11022]=47;
sine[11023]=47;
sine[11024]=47;
sine[11025]=47;
sine[11026]=47;
sine[11027]=47;
sine[11028]=47;
sine[11029]=47;
sine[11030]=47;
sine[11031]=47;
sine[11032]=47;
sine[11033]=47;
sine[11034]=47;
sine[11035]=47;
sine[11036]=47;
sine[11037]=47;
sine[11038]=47;
sine[11039]=47;
sine[11040]=47;
sine[11041]=48;
sine[11042]=48;
sine[11043]=48;
sine[11044]=48;
sine[11045]=48;
sine[11046]=48;
sine[11047]=48;
sine[11048]=48;
sine[11049]=48;
sine[11050]=48;
sine[11051]=48;
sine[11052]=48;
sine[11053]=48;
sine[11054]=48;
sine[11055]=48;
sine[11056]=48;
sine[11057]=48;
sine[11058]=48;
sine[11059]=48;
sine[11060]=48;
sine[11061]=48;
sine[11062]=48;
sine[11063]=48;
sine[11064]=48;
sine[11065]=48;
sine[11066]=49;
sine[11067]=49;
sine[11068]=49;
sine[11069]=49;
sine[11070]=49;
sine[11071]=49;
sine[11072]=49;
sine[11073]=49;
sine[11074]=49;
sine[11075]=49;
sine[11076]=49;
sine[11077]=49;
sine[11078]=49;
sine[11079]=49;
sine[11080]=49;
sine[11081]=49;
sine[11082]=49;
sine[11083]=49;
sine[11084]=49;
sine[11085]=49;
sine[11086]=49;
sine[11087]=49;
sine[11088]=49;
sine[11089]=49;
sine[11090]=49;
sine[11091]=49;
sine[11092]=49;
sine[11093]=50;
sine[11094]=50;
sine[11095]=50;
sine[11096]=50;
sine[11097]=50;
sine[11098]=50;
sine[11099]=50;
sine[11100]=50;
sine[11101]=50;
sine[11102]=50;
sine[11103]=50;
sine[11104]=50;
sine[11105]=50;
sine[11106]=50;
sine[11107]=50;
sine[11108]=50;
sine[11109]=50;
sine[11110]=50;
sine[11111]=50;
sine[11112]=50;
sine[11113]=50;
sine[11114]=50;
sine[11115]=50;
sine[11116]=50;
sine[11117]=50;
sine[11118]=50;
sine[11119]=51;
sine[11120]=51;
sine[11121]=51;
sine[11122]=51;
sine[11123]=51;
sine[11124]=51;
sine[11125]=51;
sine[11126]=51;
sine[11127]=51;
sine[11128]=51;
sine[11129]=51;
sine[11130]=51;
sine[11131]=51;
sine[11132]=51;
sine[11133]=51;
sine[11134]=51;
sine[11135]=51;
sine[11136]=51;
sine[11137]=51;
sine[11138]=51;
sine[11139]=51;
sine[11140]=51;
sine[11141]=51;
sine[11142]=51;
sine[11143]=51;
sine[11144]=51;
sine[11145]=51;
sine[11146]=52;
sine[11147]=52;
sine[11148]=52;
sine[11149]=52;
sine[11150]=52;
sine[11151]=52;
sine[11152]=52;
sine[11153]=52;
sine[11154]=52;
sine[11155]=52;
sine[11156]=52;
sine[11157]=52;
sine[11158]=52;
sine[11159]=52;
sine[11160]=52;
sine[11161]=52;
sine[11162]=52;
sine[11163]=52;
sine[11164]=52;
sine[11165]=52;
sine[11166]=52;
sine[11167]=52;
sine[11168]=52;
sine[11169]=52;
sine[11170]=52;
sine[11171]=52;
sine[11172]=52;
sine[11173]=53;
sine[11174]=53;
sine[11175]=53;
sine[11176]=53;
sine[11177]=53;
sine[11178]=53;
sine[11179]=53;
sine[11180]=53;
sine[11181]=53;
sine[11182]=53;
sine[11183]=53;
sine[11184]=53;
sine[11185]=53;
sine[11186]=53;
sine[11187]=53;
sine[11188]=53;
sine[11189]=53;
sine[11190]=53;
sine[11191]=53;
sine[11192]=53;
sine[11193]=53;
sine[11194]=53;
sine[11195]=53;
sine[11196]=53;
sine[11197]=53;
sine[11198]=53;
sine[11199]=53;
sine[11200]=53;
sine[11201]=54;
sine[11202]=54;
sine[11203]=54;
sine[11204]=54;
sine[11205]=54;
sine[11206]=54;
sine[11207]=54;
sine[11208]=54;
sine[11209]=54;
sine[11210]=54;
sine[11211]=54;
sine[11212]=54;
sine[11213]=54;
sine[11214]=54;
sine[11215]=54;
sine[11216]=54;
sine[11217]=54;
sine[11218]=54;
sine[11219]=54;
sine[11220]=54;
sine[11221]=54;
sine[11222]=54;
sine[11223]=54;
sine[11224]=54;
sine[11225]=54;
sine[11226]=54;
sine[11227]=54;
sine[11228]=54;
sine[11229]=55;
sine[11230]=55;
sine[11231]=55;
sine[11232]=55;
sine[11233]=55;
sine[11234]=55;
sine[11235]=55;
sine[11236]=55;
sine[11237]=55;
sine[11238]=55;
sine[11239]=55;
sine[11240]=55;
sine[11241]=55;
sine[11242]=55;
sine[11243]=55;
sine[11244]=55;
sine[11245]=55;
sine[11246]=55;
sine[11247]=55;
sine[11248]=55;
sine[11249]=55;
sine[11250]=55;
sine[11251]=55;
sine[11252]=55;
sine[11253]=55;
sine[11254]=55;
sine[11255]=55;
sine[11256]=55;
sine[11257]=55;
sine[11258]=56;
sine[11259]=56;
sine[11260]=56;
sine[11261]=56;
sine[11262]=56;
sine[11263]=56;
sine[11264]=56;
sine[11265]=56;
sine[11266]=56;
sine[11267]=56;
sine[11268]=56;
sine[11269]=56;
sine[11270]=56;
sine[11271]=56;
sine[11272]=56;
sine[11273]=56;
sine[11274]=56;
sine[11275]=56;
sine[11276]=56;
sine[11277]=56;
sine[11278]=56;
sine[11279]=56;
sine[11280]=56;
sine[11281]=56;
sine[11282]=56;
sine[11283]=56;
sine[11284]=56;
sine[11285]=56;
sine[11286]=56;
sine[11287]=57;
sine[11288]=57;
sine[11289]=57;
sine[11290]=57;
sine[11291]=57;
sine[11292]=57;
sine[11293]=57;
sine[11294]=57;
sine[11295]=57;
sine[11296]=57;
sine[11297]=57;
sine[11298]=57;
sine[11299]=57;
sine[11300]=57;
sine[11301]=57;
sine[11302]=57;
sine[11303]=57;
sine[11304]=57;
sine[11305]=57;
sine[11306]=57;
sine[11307]=57;
sine[11308]=57;
sine[11309]=57;
sine[11310]=57;
sine[11311]=57;
sine[11312]=57;
sine[11313]=57;
sine[11314]=57;
sine[11315]=57;
sine[11316]=57;
sine[11317]=58;
sine[11318]=58;
sine[11319]=58;
sine[11320]=58;
sine[11321]=58;
sine[11322]=58;
sine[11323]=58;
sine[11324]=58;
sine[11325]=58;
sine[11326]=58;
sine[11327]=58;
sine[11328]=58;
sine[11329]=58;
sine[11330]=58;
sine[11331]=58;
sine[11332]=58;
sine[11333]=58;
sine[11334]=58;
sine[11335]=58;
sine[11336]=58;
sine[11337]=58;
sine[11338]=58;
sine[11339]=58;
sine[11340]=58;
sine[11341]=58;
sine[11342]=58;
sine[11343]=58;
sine[11344]=58;
sine[11345]=58;
sine[11346]=58;
sine[11347]=59;
sine[11348]=59;
sine[11349]=59;
sine[11350]=59;
sine[11351]=59;
sine[11352]=59;
sine[11353]=59;
sine[11354]=59;
sine[11355]=59;
sine[11356]=59;
sine[11357]=59;
sine[11358]=59;
sine[11359]=59;
sine[11360]=59;
sine[11361]=59;
sine[11362]=59;
sine[11363]=59;
sine[11364]=59;
sine[11365]=59;
sine[11366]=59;
sine[11367]=59;
sine[11368]=59;
sine[11369]=59;
sine[11370]=59;
sine[11371]=59;
sine[11372]=59;
sine[11373]=59;
sine[11374]=59;
sine[11375]=59;
sine[11376]=59;
sine[11377]=59;
sine[11378]=60;
sine[11379]=60;
sine[11380]=60;
sine[11381]=60;
sine[11382]=60;
sine[11383]=60;
sine[11384]=60;
sine[11385]=60;
sine[11386]=60;
sine[11387]=60;
sine[11388]=60;
sine[11389]=60;
sine[11390]=60;
sine[11391]=60;
sine[11392]=60;
sine[11393]=60;
sine[11394]=60;
sine[11395]=60;
sine[11396]=60;
sine[11397]=60;
sine[11398]=60;
sine[11399]=60;
sine[11400]=60;
sine[11401]=60;
sine[11402]=60;
sine[11403]=60;
sine[11404]=60;
sine[11405]=60;
sine[11406]=60;
sine[11407]=60;
sine[11408]=60;
sine[11409]=60;
sine[11410]=61;
sine[11411]=61;
sine[11412]=61;
sine[11413]=61;
sine[11414]=61;
sine[11415]=61;
sine[11416]=61;
sine[11417]=61;
sine[11418]=61;
sine[11419]=61;
sine[11420]=61;
sine[11421]=61;
sine[11422]=61;
sine[11423]=61;
sine[11424]=61;
sine[11425]=61;
sine[11426]=61;
sine[11427]=61;
sine[11428]=61;
sine[11429]=61;
sine[11430]=61;
sine[11431]=61;
sine[11432]=61;
sine[11433]=61;
sine[11434]=61;
sine[11435]=61;
sine[11436]=61;
sine[11437]=61;
sine[11438]=61;
sine[11439]=61;
sine[11440]=61;
sine[11441]=61;
sine[11442]=61;
sine[11443]=62;
sine[11444]=62;
sine[11445]=62;
sine[11446]=62;
sine[11447]=62;
sine[11448]=62;
sine[11449]=62;
sine[11450]=62;
sine[11451]=62;
sine[11452]=62;
sine[11453]=62;
sine[11454]=62;
sine[11455]=62;
sine[11456]=62;
sine[11457]=62;
sine[11458]=62;
sine[11459]=62;
sine[11460]=62;
sine[11461]=62;
sine[11462]=62;
sine[11463]=62;
sine[11464]=62;
sine[11465]=62;
sine[11466]=62;
sine[11467]=62;
sine[11468]=62;
sine[11469]=62;
sine[11470]=62;
sine[11471]=62;
sine[11472]=62;
sine[11473]=62;
sine[11474]=62;
sine[11475]=62;
sine[11476]=63;
sine[11477]=63;
sine[11478]=63;
sine[11479]=63;
sine[11480]=63;
sine[11481]=63;
sine[11482]=63;
sine[11483]=63;
sine[11484]=63;
sine[11485]=63;
sine[11486]=63;
sine[11487]=63;
sine[11488]=63;
sine[11489]=63;
sine[11490]=63;
sine[11491]=63;
sine[11492]=63;
sine[11493]=63;
sine[11494]=63;
sine[11495]=63;
sine[11496]=63;
sine[11497]=63;
sine[11498]=63;
sine[11499]=63;
sine[11500]=63;
sine[11501]=63;
sine[11502]=63;
sine[11503]=63;
sine[11504]=63;
sine[11505]=63;
sine[11506]=63;
sine[11507]=63;
sine[11508]=63;
sine[11509]=63;
sine[11510]=63;
sine[11511]=64;
sine[11512]=64;
sine[11513]=64;
sine[11514]=64;
sine[11515]=64;
sine[11516]=64;
sine[11517]=64;
sine[11518]=64;
sine[11519]=64;
sine[11520]=64;
sine[11521]=64;
sine[11522]=64;
sine[11523]=64;
sine[11524]=64;
sine[11525]=64;
sine[11526]=64;
sine[11527]=64;
sine[11528]=64;
sine[11529]=64;
sine[11530]=64;
sine[11531]=64;
sine[11532]=64;
sine[11533]=64;
sine[11534]=64;
sine[11535]=64;
sine[11536]=64;
sine[11537]=64;
sine[11538]=64;
sine[11539]=64;
sine[11540]=64;
sine[11541]=64;
sine[11542]=64;
sine[11543]=64;
sine[11544]=64;
sine[11545]=64;
sine[11546]=65;
sine[11547]=65;
sine[11548]=65;
sine[11549]=65;
sine[11550]=65;
sine[11551]=65;
sine[11552]=65;
sine[11553]=65;
sine[11554]=65;
sine[11555]=65;
sine[11556]=65;
sine[11557]=65;
sine[11558]=65;
sine[11559]=65;
sine[11560]=65;
sine[11561]=65;
sine[11562]=65;
sine[11563]=65;
sine[11564]=65;
sine[11565]=65;
sine[11566]=65;
sine[11567]=65;
sine[11568]=65;
sine[11569]=65;
sine[11570]=65;
sine[11571]=65;
sine[11572]=65;
sine[11573]=65;
sine[11574]=65;
sine[11575]=65;
sine[11576]=65;
sine[11577]=65;
sine[11578]=65;
sine[11579]=65;
sine[11580]=65;
sine[11581]=65;
sine[11582]=65;
sine[11583]=66;
sine[11584]=66;
sine[11585]=66;
sine[11586]=66;
sine[11587]=66;
sine[11588]=66;
sine[11589]=66;
sine[11590]=66;
sine[11591]=66;
sine[11592]=66;
sine[11593]=66;
sine[11594]=66;
sine[11595]=66;
sine[11596]=66;
sine[11597]=66;
sine[11598]=66;
sine[11599]=66;
sine[11600]=66;
sine[11601]=66;
sine[11602]=66;
sine[11603]=66;
sine[11604]=66;
sine[11605]=66;
sine[11606]=66;
sine[11607]=66;
sine[11608]=66;
sine[11609]=66;
sine[11610]=66;
sine[11611]=66;
sine[11612]=66;
sine[11613]=66;
sine[11614]=66;
sine[11615]=66;
sine[11616]=66;
sine[11617]=66;
sine[11618]=66;
sine[11619]=66;
sine[11620]=66;
sine[11621]=67;
sine[11622]=67;
sine[11623]=67;
sine[11624]=67;
sine[11625]=67;
sine[11626]=67;
sine[11627]=67;
sine[11628]=67;
sine[11629]=67;
sine[11630]=67;
sine[11631]=67;
sine[11632]=67;
sine[11633]=67;
sine[11634]=67;
sine[11635]=67;
sine[11636]=67;
sine[11637]=67;
sine[11638]=67;
sine[11639]=67;
sine[11640]=67;
sine[11641]=67;
sine[11642]=67;
sine[11643]=67;
sine[11644]=67;
sine[11645]=67;
sine[11646]=67;
sine[11647]=67;
sine[11648]=67;
sine[11649]=67;
sine[11650]=67;
sine[11651]=67;
sine[11652]=67;
sine[11653]=67;
sine[11654]=67;
sine[11655]=67;
sine[11656]=67;
sine[11657]=67;
sine[11658]=67;
sine[11659]=67;
sine[11660]=67;
sine[11661]=68;
sine[11662]=68;
sine[11663]=68;
sine[11664]=68;
sine[11665]=68;
sine[11666]=68;
sine[11667]=68;
sine[11668]=68;
sine[11669]=68;
sine[11670]=68;
sine[11671]=68;
sine[11672]=68;
sine[11673]=68;
sine[11674]=68;
sine[11675]=68;
sine[11676]=68;
sine[11677]=68;
sine[11678]=68;
sine[11679]=68;
sine[11680]=68;
sine[11681]=68;
sine[11682]=68;
sine[11683]=68;
sine[11684]=68;
sine[11685]=68;
sine[11686]=68;
sine[11687]=68;
sine[11688]=68;
sine[11689]=68;
sine[11690]=68;
sine[11691]=68;
sine[11692]=68;
sine[11693]=68;
sine[11694]=68;
sine[11695]=68;
sine[11696]=68;
sine[11697]=68;
sine[11698]=68;
sine[11699]=68;
sine[11700]=68;
sine[11701]=68;
sine[11702]=69;
sine[11703]=69;
sine[11704]=69;
sine[11705]=69;
sine[11706]=69;
sine[11707]=69;
sine[11708]=69;
sine[11709]=69;
sine[11710]=69;
sine[11711]=69;
sine[11712]=69;
sine[11713]=69;
sine[11714]=69;
sine[11715]=69;
sine[11716]=69;
sine[11717]=69;
sine[11718]=69;
sine[11719]=69;
sine[11720]=69;
sine[11721]=69;
sine[11722]=69;
sine[11723]=69;
sine[11724]=69;
sine[11725]=69;
sine[11726]=69;
sine[11727]=69;
sine[11728]=69;
sine[11729]=69;
sine[11730]=69;
sine[11731]=69;
sine[11732]=69;
sine[11733]=69;
sine[11734]=69;
sine[11735]=69;
sine[11736]=69;
sine[11737]=69;
sine[11738]=69;
sine[11739]=69;
sine[11740]=69;
sine[11741]=69;
sine[11742]=69;
sine[11743]=69;
sine[11744]=69;
sine[11745]=69;
sine[11746]=70;
sine[11747]=70;
sine[11748]=70;
sine[11749]=70;
sine[11750]=70;
sine[11751]=70;
sine[11752]=70;
sine[11753]=70;
sine[11754]=70;
sine[11755]=70;
sine[11756]=70;
sine[11757]=70;
sine[11758]=70;
sine[11759]=70;
sine[11760]=70;
sine[11761]=70;
sine[11762]=70;
sine[11763]=70;
sine[11764]=70;
sine[11765]=70;
sine[11766]=70;
sine[11767]=70;
sine[11768]=70;
sine[11769]=70;
sine[11770]=70;
sine[11771]=70;
sine[11772]=70;
sine[11773]=70;
sine[11774]=70;
sine[11775]=70;
sine[11776]=70;
sine[11777]=70;
sine[11778]=70;
sine[11779]=70;
sine[11780]=70;
sine[11781]=70;
sine[11782]=70;
sine[11783]=70;
sine[11784]=70;
sine[11785]=70;
sine[11786]=70;
sine[11787]=70;
sine[11788]=70;
sine[11789]=70;
sine[11790]=70;
sine[11791]=71;
sine[11792]=71;
sine[11793]=71;
sine[11794]=71;
sine[11795]=71;
sine[11796]=71;
sine[11797]=71;
sine[11798]=71;
sine[11799]=71;
sine[11800]=71;
sine[11801]=71;
sine[11802]=71;
sine[11803]=71;
sine[11804]=71;
sine[11805]=71;
sine[11806]=71;
sine[11807]=71;
sine[11808]=71;
sine[11809]=71;
sine[11810]=71;
sine[11811]=71;
sine[11812]=71;
sine[11813]=71;
sine[11814]=71;
sine[11815]=71;
sine[11816]=71;
sine[11817]=71;
sine[11818]=71;
sine[11819]=71;
sine[11820]=71;
sine[11821]=71;
sine[11822]=71;
sine[11823]=71;
sine[11824]=71;
sine[11825]=71;
sine[11826]=71;
sine[11827]=71;
sine[11828]=71;
sine[11829]=71;
sine[11830]=71;
sine[11831]=71;
sine[11832]=71;
sine[11833]=71;
sine[11834]=71;
sine[11835]=71;
sine[11836]=71;
sine[11837]=71;
sine[11838]=71;
sine[11839]=71;
sine[11840]=72;
sine[11841]=72;
sine[11842]=72;
sine[11843]=72;
sine[11844]=72;
sine[11845]=72;
sine[11846]=72;
sine[11847]=72;
sine[11848]=72;
sine[11849]=72;
sine[11850]=72;
sine[11851]=72;
sine[11852]=72;
sine[11853]=72;
sine[11854]=72;
sine[11855]=72;
sine[11856]=72;
sine[11857]=72;
sine[11858]=72;
sine[11859]=72;
sine[11860]=72;
sine[11861]=72;
sine[11862]=72;
sine[11863]=72;
sine[11864]=72;
sine[11865]=72;
sine[11866]=72;
sine[11867]=72;
sine[11868]=72;
sine[11869]=72;
sine[11870]=72;
sine[11871]=72;
sine[11872]=72;
sine[11873]=72;
sine[11874]=72;
sine[11875]=72;
sine[11876]=72;
sine[11877]=72;
sine[11878]=72;
sine[11879]=72;
sine[11880]=72;
sine[11881]=72;
sine[11882]=72;
sine[11883]=72;
sine[11884]=72;
sine[11885]=72;
sine[11886]=72;
sine[11887]=72;
sine[11888]=72;
sine[11889]=72;
sine[11890]=72;
sine[11891]=72;
sine[11892]=72;
sine[11893]=73;
sine[11894]=73;
sine[11895]=73;
sine[11896]=73;
sine[11897]=73;
sine[11898]=73;
sine[11899]=73;
sine[11900]=73;
sine[11901]=73;
sine[11902]=73;
sine[11903]=73;
sine[11904]=73;
sine[11905]=73;
sine[11906]=73;
sine[11907]=73;
sine[11908]=73;
sine[11909]=73;
sine[11910]=73;
sine[11911]=73;
sine[11912]=73;
sine[11913]=73;
sine[11914]=73;
sine[11915]=73;
sine[11916]=73;
sine[11917]=73;
sine[11918]=73;
sine[11919]=73;
sine[11920]=73;
sine[11921]=73;
sine[11922]=73;
sine[11923]=73;
sine[11924]=73;
sine[11925]=73;
sine[11926]=73;
sine[11927]=73;
sine[11928]=73;
sine[11929]=73;
sine[11930]=73;
sine[11931]=73;
sine[11932]=73;
sine[11933]=73;
sine[11934]=73;
sine[11935]=73;
sine[11936]=73;
sine[11937]=73;
sine[11938]=73;
sine[11939]=73;
sine[11940]=73;
sine[11941]=73;
sine[11942]=73;
sine[11943]=73;
sine[11944]=73;
sine[11945]=73;
sine[11946]=73;
sine[11947]=73;
sine[11948]=73;
sine[11949]=73;
sine[11950]=74;
sine[11951]=74;
sine[11952]=74;
sine[11953]=74;
sine[11954]=74;
sine[11955]=74;
sine[11956]=74;
sine[11957]=74;
sine[11958]=74;
sine[11959]=74;
sine[11960]=74;
sine[11961]=74;
sine[11962]=74;
sine[11963]=74;
sine[11964]=74;
sine[11965]=74;
sine[11966]=74;
sine[11967]=74;
sine[11968]=74;
sine[11969]=74;
sine[11970]=74;
sine[11971]=74;
sine[11972]=74;
sine[11973]=74;
sine[11974]=74;
sine[11975]=74;
sine[11976]=74;
sine[11977]=74;
sine[11978]=74;
sine[11979]=74;
sine[11980]=74;
sine[11981]=74;
sine[11982]=74;
sine[11983]=74;
sine[11984]=74;
sine[11985]=74;
sine[11986]=74;
sine[11987]=74;
sine[11988]=74;
sine[11989]=74;
sine[11990]=74;
sine[11991]=74;
sine[11992]=74;
sine[11993]=74;
sine[11994]=74;
sine[11995]=74;
sine[11996]=74;
sine[11997]=74;
sine[11998]=74;
sine[11999]=74;
sine[12000]=74;
sine[12001]=74;
sine[12002]=74;
sine[12003]=74;
sine[12004]=74;
sine[12005]=74;
sine[12006]=74;
sine[12007]=74;
sine[12008]=74;
sine[12009]=74;
sine[12010]=74;
sine[12011]=74;
sine[12012]=74;
sine[12013]=74;
sine[12014]=75;
sine[12015]=75;
sine[12016]=75;
sine[12017]=75;
sine[12018]=75;
sine[12019]=75;
sine[12020]=75;
sine[12021]=75;
sine[12022]=75;
sine[12023]=75;
sine[12024]=75;
sine[12025]=75;
sine[12026]=75;
sine[12027]=75;
sine[12028]=75;
sine[12029]=75;
sine[12030]=75;
sine[12031]=75;
sine[12032]=75;
sine[12033]=75;
sine[12034]=75;
sine[12035]=75;
sine[12036]=75;
sine[12037]=75;
sine[12038]=75;
sine[12039]=75;
sine[12040]=75;
sine[12041]=75;
sine[12042]=75;
sine[12043]=75;
sine[12044]=75;
sine[12045]=75;
sine[12046]=75;
sine[12047]=75;
sine[12048]=75;
sine[12049]=75;
sine[12050]=75;
sine[12051]=75;
sine[12052]=75;
sine[12053]=75;
sine[12054]=75;
sine[12055]=75;
sine[12056]=75;
sine[12057]=75;
sine[12058]=75;
sine[12059]=75;
sine[12060]=75;
sine[12061]=75;
sine[12062]=75;
sine[12063]=75;
sine[12064]=75;
sine[12065]=75;
sine[12066]=75;
sine[12067]=75;
sine[12068]=75;
sine[12069]=75;
sine[12070]=75;
sine[12071]=75;
sine[12072]=75;
sine[12073]=75;
sine[12074]=75;
sine[12075]=75;
sine[12076]=75;
sine[12077]=75;
sine[12078]=75;
sine[12079]=75;
sine[12080]=75;
sine[12081]=75;
sine[12082]=75;
sine[12083]=75;
sine[12084]=75;
sine[12085]=75;
sine[12086]=75;
sine[12087]=76;
sine[12088]=76;
sine[12089]=76;
sine[12090]=76;
sine[12091]=76;
sine[12092]=76;
sine[12093]=76;
sine[12094]=76;
sine[12095]=76;
sine[12096]=76;
sine[12097]=76;
sine[12098]=76;
sine[12099]=76;
sine[12100]=76;
sine[12101]=76;
sine[12102]=76;
sine[12103]=76;
sine[12104]=76;
sine[12105]=76;
sine[12106]=76;
sine[12107]=76;
sine[12108]=76;
sine[12109]=76;
sine[12110]=76;
sine[12111]=76;
sine[12112]=76;
sine[12113]=76;
sine[12114]=76;
sine[12115]=76;
sine[12116]=76;
sine[12117]=76;
sine[12118]=76;
sine[12119]=76;
sine[12120]=76;
sine[12121]=76;
sine[12122]=76;
sine[12123]=76;
sine[12124]=76;
sine[12125]=76;
sine[12126]=76;
sine[12127]=76;
sine[12128]=76;
sine[12129]=76;
sine[12130]=76;
sine[12131]=76;
sine[12132]=76;
sine[12133]=76;
sine[12134]=76;
sine[12135]=76;
sine[12136]=76;
sine[12137]=76;
sine[12138]=76;
sine[12139]=76;
sine[12140]=76;
sine[12141]=76;
sine[12142]=76;
sine[12143]=76;
sine[12144]=76;
sine[12145]=76;
sine[12146]=76;
sine[12147]=76;
sine[12148]=76;
sine[12149]=76;
sine[12150]=76;
sine[12151]=76;
sine[12152]=76;
sine[12153]=76;
sine[12154]=76;
sine[12155]=76;
sine[12156]=76;
sine[12157]=76;
sine[12158]=76;
sine[12159]=76;
sine[12160]=76;
sine[12161]=76;
sine[12162]=76;
sine[12163]=76;
sine[12164]=76;
sine[12165]=76;
sine[12166]=76;
sine[12167]=76;
sine[12168]=76;
sine[12169]=76;
sine[12170]=76;
sine[12171]=76;
sine[12172]=76;
sine[12173]=76;
sine[12174]=76;
sine[12175]=77;
sine[12176]=77;
sine[12177]=77;
sine[12178]=77;
sine[12179]=77;
sine[12180]=77;
sine[12181]=77;
sine[12182]=77;
sine[12183]=77;
sine[12184]=77;
sine[12185]=77;
sine[12186]=77;
sine[12187]=77;
sine[12188]=77;
sine[12189]=77;
sine[12190]=77;
sine[12191]=77;
sine[12192]=77;
sine[12193]=77;
sine[12194]=77;
sine[12195]=77;
sine[12196]=77;
sine[12197]=77;
sine[12198]=77;
sine[12199]=77;
sine[12200]=77;
sine[12201]=77;
sine[12202]=77;
sine[12203]=77;
sine[12204]=77;
sine[12205]=77;
sine[12206]=77;
sine[12207]=77;
sine[12208]=77;
sine[12209]=77;
sine[12210]=77;
sine[12211]=77;
sine[12212]=77;
sine[12213]=77;
sine[12214]=77;
sine[12215]=77;
sine[12216]=77;
sine[12217]=77;
sine[12218]=77;
sine[12219]=77;
sine[12220]=77;
sine[12221]=77;
sine[12222]=77;
sine[12223]=77;
sine[12224]=77;
sine[12225]=77;
sine[12226]=77;
sine[12227]=77;
sine[12228]=77;
sine[12229]=77;
sine[12230]=77;
sine[12231]=77;
sine[12232]=77;
sine[12233]=77;
sine[12234]=77;
sine[12235]=77;
sine[12236]=77;
sine[12237]=77;
sine[12238]=77;
sine[12239]=77;
sine[12240]=77;
sine[12241]=77;
sine[12242]=77;
sine[12243]=77;
sine[12244]=77;
sine[12245]=77;
sine[12246]=77;
sine[12247]=77;
sine[12248]=77;
sine[12249]=77;
sine[12250]=77;
sine[12251]=77;
sine[12252]=77;
sine[12253]=77;
sine[12254]=77;
sine[12255]=77;
sine[12256]=77;
sine[12257]=77;
sine[12258]=77;
sine[12259]=77;
sine[12260]=77;
sine[12261]=77;
sine[12262]=77;
sine[12263]=77;
sine[12264]=77;
sine[12265]=77;
sine[12266]=77;
sine[12267]=77;
sine[12268]=77;
sine[12269]=77;
sine[12270]=77;
sine[12271]=77;
sine[12272]=77;
sine[12273]=77;
sine[12274]=77;
sine[12275]=77;
sine[12276]=77;
sine[12277]=77;
sine[12278]=77;
sine[12279]=77;
sine[12280]=77;
sine[12281]=77;
sine[12282]=77;
sine[12283]=77;
sine[12284]=77;
sine[12285]=77;
sine[12286]=77;
sine[12287]=77;
sine[12288]=77;
sine[12289]=77;
sine[12290]=77;
sine[12291]=77;
sine[12292]=77;
sine[12293]=77;
sine[12294]=77;
sine[12295]=77;
sine[12296]=77;
sine[12297]=77;
sine[12298]=77;
sine[12299]=78;
sine[12300]=78;
sine[12301]=78;
sine[12302]=78;
sine[12303]=78;
sine[12304]=78;
sine[12305]=78;
sine[12306]=78;
sine[12307]=78;
sine[12308]=78;
sine[12309]=78;
sine[12310]=78;
sine[12311]=78;
sine[12312]=78;
sine[12313]=78;
sine[12314]=78;
sine[12315]=78;
sine[12316]=78;
sine[12317]=78;
sine[12318]=78;
sine[12319]=78;
sine[12320]=78;
sine[12321]=78;
sine[12322]=78;
sine[12323]=78;
sine[12324]=78;
sine[12325]=78;
sine[12326]=78;
sine[12327]=78;
sine[12328]=78;
sine[12329]=78;
sine[12330]=78;
sine[12331]=78;
sine[12332]=78;
sine[12333]=78;
sine[12334]=78;
sine[12335]=78;
sine[12336]=78;
sine[12337]=78;
sine[12338]=78;
sine[12339]=78;
sine[12340]=78;
sine[12341]=78;
sine[12342]=78;
sine[12343]=78;
sine[12344]=78;
sine[12345]=78;
sine[12346]=78;
sine[12347]=78;
sine[12348]=78;
sine[12349]=78;
sine[12350]=78;
sine[12351]=78;
sine[12352]=78;
sine[12353]=78;
sine[12354]=78;
sine[12355]=78;
sine[12356]=78;
sine[12357]=78;
sine[12358]=78;
sine[12359]=78;
sine[12360]=78;
sine[12361]=78;
sine[12362]=78;
sine[12363]=78;
sine[12364]=78;
sine[12365]=78;
sine[12366]=78;
sine[12367]=78;
sine[12368]=78;
sine[12369]=78;
sine[12370]=78;
sine[12371]=78;
sine[12372]=78;
sine[12373]=78;
sine[12374]=78;
sine[12375]=78;
sine[12376]=78;
sine[12377]=78;
sine[12378]=78;
sine[12379]=78;
sine[12380]=78;
sine[12381]=78;
sine[12382]=78;
sine[12383]=78;
sine[12384]=78;
sine[12385]=78;
sine[12386]=78;
sine[12387]=78;
sine[12388]=78;
sine[12389]=78;
sine[12390]=78;
sine[12391]=78;
sine[12392]=78;
sine[12393]=78;
sine[12394]=78;
sine[12395]=78;
sine[12396]=78;
sine[12397]=78;
sine[12398]=78;
sine[12399]=78;
sine[12400]=78;
sine[12401]=78;
sine[12402]=78;
sine[12403]=78;
sine[12404]=78;
sine[12405]=78;
sine[12406]=78;
sine[12407]=78;
sine[12408]=78;
sine[12409]=78;
sine[12410]=78;
sine[12411]=78;
sine[12412]=78;
sine[12413]=78;
sine[12414]=78;
sine[12415]=78;
sine[12416]=78;
sine[12417]=78;
sine[12418]=78;
sine[12419]=78;
sine[12420]=78;
sine[12421]=78;
sine[12422]=78;
sine[12423]=78;
sine[12424]=78;
sine[12425]=78;
sine[12426]=78;
sine[12427]=78;
sine[12428]=78;
sine[12429]=78;
sine[12430]=78;
sine[12431]=78;
sine[12432]=78;
sine[12433]=78;
sine[12434]=78;
sine[12435]=78;
sine[12436]=78;
sine[12437]=78;
sine[12438]=78;
sine[12439]=78;
sine[12440]=78;
sine[12441]=78;
sine[12442]=78;
sine[12443]=78;
sine[12444]=78;
sine[12445]=78;
sine[12446]=78;
sine[12447]=78;
sine[12448]=78;
sine[12449]=78;
sine[12450]=78;
sine[12451]=78;
sine[12452]=78;
sine[12453]=78;
sine[12454]=78;
sine[12455]=78;
sine[12456]=78;
sine[12457]=78;
sine[12458]=78;
sine[12459]=78;
sine[12460]=78;
sine[12461]=78;
sine[12462]=78;
sine[12463]=78;
sine[12464]=78;
sine[12465]=78;
sine[12466]=78;
sine[12467]=78;
sine[12468]=78;
sine[12469]=78;
sine[12470]=78;
sine[12471]=78;
sine[12472]=78;
sine[12473]=78;
sine[12474]=78;
sine[12475]=78;
sine[12476]=78;
sine[12477]=78;
sine[12478]=78;
sine[12479]=78;
sine[12480]=78;
sine[12481]=78;
sine[12482]=78;
sine[12483]=78;
sine[12484]=78;
sine[12485]=78;
sine[12486]=78;
sine[12487]=78;
sine[12488]=78;
sine[12489]=78;
sine[12490]=78;
sine[12491]=78;
sine[12492]=78;
sine[12493]=78;
sine[12494]=78;
sine[12495]=78;
sine[12496]=78;
sine[12497]=78;
sine[12498]=78;
sine[12499]=78;
sine[12500]=78;
sine[12501]=78;
sine[12502]=78;
sine[12503]=78;
sine[12504]=78;
sine[12505]=78;
sine[12506]=78;
sine[12507]=78;
sine[12508]=78;
sine[12509]=78;
sine[12510]=78;
sine[12511]=78;
sine[12512]=78;
sine[12513]=78;
sine[12514]=78;
sine[12515]=78;
sine[12516]=78;
sine[12517]=78;
sine[12518]=78;
sine[12519]=78;
sine[12520]=78;
sine[12521]=78;
sine[12522]=78;
sine[12523]=78;
sine[12524]=78;
sine[12525]=78;
sine[12526]=78;
sine[12527]=78;
sine[12528]=78;
sine[12529]=78;
sine[12530]=78;
sine[12531]=78;
sine[12532]=78;
sine[12533]=78;
sine[12534]=78;
sine[12535]=78;
sine[12536]=78;
sine[12537]=78;
sine[12538]=78;
sine[12539]=78;
sine[12540]=78;
sine[12541]=78;
sine[12542]=78;
sine[12543]=78;
sine[12544]=78;
sine[12545]=78;
sine[12546]=78;
sine[12547]=78;
sine[12548]=78;
sine[12549]=78;
sine[12550]=78;
sine[12551]=78;
sine[12552]=78;
sine[12553]=78;
sine[12554]=78;
sine[12555]=78;
sine[12556]=78;
sine[12557]=78;
sine[12558]=78;
sine[12559]=78;
sine[12560]=78;
sine[12561]=78;
sine[12562]=78;
sine[12563]=78;
sine[12564]=78;
sine[12565]=78;
sine[12566]=78;
sine[12567]=78;
sine[12568]=78;
sine[12569]=78;
sine[12570]=78;
sine[12571]=78;
sine[12572]=78;
sine[12573]=78;
sine[12574]=78;
sine[12575]=78;
sine[12576]=78;
sine[12577]=78;
sine[12578]=78;
sine[12579]=78;
sine[12580]=78;
sine[12581]=78;
sine[12582]=78;
sine[12583]=78;
sine[12584]=78;
sine[12585]=78;
sine[12586]=78;
sine[12587]=78;
sine[12588]=78;
sine[12589]=78;
sine[12590]=78;
sine[12591]=78;
sine[12592]=78;
sine[12593]=78;
sine[12594]=78;
sine[12595]=78;
sine[12596]=78;
sine[12597]=78;
sine[12598]=78;
sine[12599]=78;
sine[12600]=78;
sine[12601]=78;
sine[12602]=78;
sine[12603]=78;
sine[12604]=78;
sine[12605]=78;
sine[12606]=78;
sine[12607]=78;
sine[12608]=78;
sine[12609]=78;
sine[12610]=78;
sine[12611]=78;
sine[12612]=78;
sine[12613]=78;
sine[12614]=78;
sine[12615]=78;
sine[12616]=78;
sine[12617]=78;
sine[12618]=78;
sine[12619]=78;
sine[12620]=78;
sine[12621]=78;
sine[12622]=78;
sine[12623]=78;
sine[12624]=78;
sine[12625]=78;
sine[12626]=78;
sine[12627]=78;
sine[12628]=78;
sine[12629]=78;
sine[12630]=78;
sine[12631]=78;
sine[12632]=78;
sine[12633]=78;
sine[12634]=78;
sine[12635]=78;
sine[12636]=78;
sine[12637]=78;
sine[12638]=78;
sine[12639]=78;
sine[12640]=78;
sine[12641]=78;
sine[12642]=78;
sine[12643]=78;
sine[12644]=78;
sine[12645]=78;
sine[12646]=78;
sine[12647]=78;
sine[12648]=78;
sine[12649]=78;
sine[12650]=78;
sine[12651]=78;
sine[12652]=78;
sine[12653]=78;
sine[12654]=78;
sine[12655]=78;
sine[12656]=78;
sine[12657]=78;
sine[12658]=78;
sine[12659]=78;
sine[12660]=78;
sine[12661]=78;
sine[12662]=78;
sine[12663]=78;
sine[12664]=78;
sine[12665]=78;
sine[12666]=78;
sine[12667]=78;
sine[12668]=78;
sine[12669]=78;
sine[12670]=78;
sine[12671]=78;
sine[12672]=78;
sine[12673]=78;
sine[12674]=78;
sine[12675]=78;
sine[12676]=78;
sine[12677]=78;
sine[12678]=78;
sine[12679]=78;
sine[12680]=78;
sine[12681]=78;
sine[12682]=78;
sine[12683]=78;
sine[12684]=78;
sine[12685]=78;
sine[12686]=78;
sine[12687]=78;
sine[12688]=78;
sine[12689]=78;
sine[12690]=78;
sine[12691]=78;
sine[12692]=78;
sine[12693]=78;
sine[12694]=78;
sine[12695]=78;
sine[12696]=78;
sine[12697]=78;
sine[12698]=78;
sine[12699]=78;
sine[12700]=78;
sine[12701]=78;
sine[12702]=77;
sine[12703]=77;
sine[12704]=77;
sine[12705]=77;
sine[12706]=77;
sine[12707]=77;
sine[12708]=77;
sine[12709]=77;
sine[12710]=77;
sine[12711]=77;
sine[12712]=77;
sine[12713]=77;
sine[12714]=77;
sine[12715]=77;
sine[12716]=77;
sine[12717]=77;
sine[12718]=77;
sine[12719]=77;
sine[12720]=77;
sine[12721]=77;
sine[12722]=77;
sine[12723]=77;
sine[12724]=77;
sine[12725]=77;
sine[12726]=77;
sine[12727]=77;
sine[12728]=77;
sine[12729]=77;
sine[12730]=77;
sine[12731]=77;
sine[12732]=77;
sine[12733]=77;
sine[12734]=77;
sine[12735]=77;
sine[12736]=77;
sine[12737]=77;
sine[12738]=77;
sine[12739]=77;
sine[12740]=77;
sine[12741]=77;
sine[12742]=77;
sine[12743]=77;
sine[12744]=77;
sine[12745]=77;
sine[12746]=77;
sine[12747]=77;
sine[12748]=77;
sine[12749]=77;
sine[12750]=77;
sine[12751]=77;
sine[12752]=77;
sine[12753]=77;
sine[12754]=77;
sine[12755]=77;
sine[12756]=77;
sine[12757]=77;
sine[12758]=77;
sine[12759]=77;
sine[12760]=77;
sine[12761]=77;
sine[12762]=77;
sine[12763]=77;
sine[12764]=77;
sine[12765]=77;
sine[12766]=77;
sine[12767]=77;
sine[12768]=77;
sine[12769]=77;
sine[12770]=77;
sine[12771]=77;
sine[12772]=77;
sine[12773]=77;
sine[12774]=77;
sine[12775]=77;
sine[12776]=77;
sine[12777]=77;
sine[12778]=77;
sine[12779]=77;
sine[12780]=77;
sine[12781]=77;
sine[12782]=77;
sine[12783]=77;
sine[12784]=77;
sine[12785]=77;
sine[12786]=77;
sine[12787]=77;
sine[12788]=77;
sine[12789]=77;
sine[12790]=77;
sine[12791]=77;
sine[12792]=77;
sine[12793]=77;
sine[12794]=77;
sine[12795]=77;
sine[12796]=77;
sine[12797]=77;
sine[12798]=77;
sine[12799]=77;
sine[12800]=77;
sine[12801]=77;
sine[12802]=77;
sine[12803]=77;
sine[12804]=77;
sine[12805]=77;
sine[12806]=77;
sine[12807]=77;
sine[12808]=77;
sine[12809]=77;
sine[12810]=77;
sine[12811]=77;
sine[12812]=77;
sine[12813]=77;
sine[12814]=77;
sine[12815]=77;
sine[12816]=77;
sine[12817]=77;
sine[12818]=77;
sine[12819]=77;
sine[12820]=77;
sine[12821]=77;
sine[12822]=77;
sine[12823]=77;
sine[12824]=77;
sine[12825]=77;
sine[12826]=76;
sine[12827]=76;
sine[12828]=76;
sine[12829]=76;
sine[12830]=76;
sine[12831]=76;
sine[12832]=76;
sine[12833]=76;
sine[12834]=76;
sine[12835]=76;
sine[12836]=76;
sine[12837]=76;
sine[12838]=76;
sine[12839]=76;
sine[12840]=76;
sine[12841]=76;
sine[12842]=76;
sine[12843]=76;
sine[12844]=76;
sine[12845]=76;
sine[12846]=76;
sine[12847]=76;
sine[12848]=76;
sine[12849]=76;
sine[12850]=76;
sine[12851]=76;
sine[12852]=76;
sine[12853]=76;
sine[12854]=76;
sine[12855]=76;
sine[12856]=76;
sine[12857]=76;
sine[12858]=76;
sine[12859]=76;
sine[12860]=76;
sine[12861]=76;
sine[12862]=76;
sine[12863]=76;
sine[12864]=76;
sine[12865]=76;
sine[12866]=76;
sine[12867]=76;
sine[12868]=76;
sine[12869]=76;
sine[12870]=76;
sine[12871]=76;
sine[12872]=76;
sine[12873]=76;
sine[12874]=76;
sine[12875]=76;
sine[12876]=76;
sine[12877]=76;
sine[12878]=76;
sine[12879]=76;
sine[12880]=76;
sine[12881]=76;
sine[12882]=76;
sine[12883]=76;
sine[12884]=76;
sine[12885]=76;
sine[12886]=76;
sine[12887]=76;
sine[12888]=76;
sine[12889]=76;
sine[12890]=76;
sine[12891]=76;
sine[12892]=76;
sine[12893]=76;
sine[12894]=76;
sine[12895]=76;
sine[12896]=76;
sine[12897]=76;
sine[12898]=76;
sine[12899]=76;
sine[12900]=76;
sine[12901]=76;
sine[12902]=76;
sine[12903]=76;
sine[12904]=76;
sine[12905]=76;
sine[12906]=76;
sine[12907]=76;
sine[12908]=76;
sine[12909]=76;
sine[12910]=76;
sine[12911]=76;
sine[12912]=76;
sine[12913]=76;
sine[12914]=75;
sine[12915]=75;
sine[12916]=75;
sine[12917]=75;
sine[12918]=75;
sine[12919]=75;
sine[12920]=75;
sine[12921]=75;
sine[12922]=75;
sine[12923]=75;
sine[12924]=75;
sine[12925]=75;
sine[12926]=75;
sine[12927]=75;
sine[12928]=75;
sine[12929]=75;
sine[12930]=75;
sine[12931]=75;
sine[12932]=75;
sine[12933]=75;
sine[12934]=75;
sine[12935]=75;
sine[12936]=75;
sine[12937]=75;
sine[12938]=75;
sine[12939]=75;
sine[12940]=75;
sine[12941]=75;
sine[12942]=75;
sine[12943]=75;
sine[12944]=75;
sine[12945]=75;
sine[12946]=75;
sine[12947]=75;
sine[12948]=75;
sine[12949]=75;
sine[12950]=75;
sine[12951]=75;
sine[12952]=75;
sine[12953]=75;
sine[12954]=75;
sine[12955]=75;
sine[12956]=75;
sine[12957]=75;
sine[12958]=75;
sine[12959]=75;
sine[12960]=75;
sine[12961]=75;
sine[12962]=75;
sine[12963]=75;
sine[12964]=75;
sine[12965]=75;
sine[12966]=75;
sine[12967]=75;
sine[12968]=75;
sine[12969]=75;
sine[12970]=75;
sine[12971]=75;
sine[12972]=75;
sine[12973]=75;
sine[12974]=75;
sine[12975]=75;
sine[12976]=75;
sine[12977]=75;
sine[12978]=75;
sine[12979]=75;
sine[12980]=75;
sine[12981]=75;
sine[12982]=75;
sine[12983]=75;
sine[12984]=75;
sine[12985]=75;
sine[12986]=75;
sine[12987]=74;
sine[12988]=74;
sine[12989]=74;
sine[12990]=74;
sine[12991]=74;
sine[12992]=74;
sine[12993]=74;
sine[12994]=74;
sine[12995]=74;
sine[12996]=74;
sine[12997]=74;
sine[12998]=74;
sine[12999]=74;
sine[13000]=74;
sine[13001]=74;
sine[13002]=74;
sine[13003]=74;
sine[13004]=74;
sine[13005]=74;
sine[13006]=74;
sine[13007]=74;
sine[13008]=74;
sine[13009]=74;
sine[13010]=74;
sine[13011]=74;
sine[13012]=74;
sine[13013]=74;
sine[13014]=74;
sine[13015]=74;
sine[13016]=74;
sine[13017]=74;
sine[13018]=74;
sine[13019]=74;
sine[13020]=74;
sine[13021]=74;
sine[13022]=74;
sine[13023]=74;
sine[13024]=74;
sine[13025]=74;
sine[13026]=74;
sine[13027]=74;
sine[13028]=74;
sine[13029]=74;
sine[13030]=74;
sine[13031]=74;
sine[13032]=74;
sine[13033]=74;
sine[13034]=74;
sine[13035]=74;
sine[13036]=74;
sine[13037]=74;
sine[13038]=74;
sine[13039]=74;
sine[13040]=74;
sine[13041]=74;
sine[13042]=74;
sine[13043]=74;
sine[13044]=74;
sine[13045]=74;
sine[13046]=74;
sine[13047]=74;
sine[13048]=74;
sine[13049]=74;
sine[13050]=74;
sine[13051]=73;
sine[13052]=73;
sine[13053]=73;
sine[13054]=73;
sine[13055]=73;
sine[13056]=73;
sine[13057]=73;
sine[13058]=73;
sine[13059]=73;
sine[13060]=73;
sine[13061]=73;
sine[13062]=73;
sine[13063]=73;
sine[13064]=73;
sine[13065]=73;
sine[13066]=73;
sine[13067]=73;
sine[13068]=73;
sine[13069]=73;
sine[13070]=73;
sine[13071]=73;
sine[13072]=73;
sine[13073]=73;
sine[13074]=73;
sine[13075]=73;
sine[13076]=73;
sine[13077]=73;
sine[13078]=73;
sine[13079]=73;
sine[13080]=73;
sine[13081]=73;
sine[13082]=73;
sine[13083]=73;
sine[13084]=73;
sine[13085]=73;
sine[13086]=73;
sine[13087]=73;
sine[13088]=73;
sine[13089]=73;
sine[13090]=73;
sine[13091]=73;
sine[13092]=73;
sine[13093]=73;
sine[13094]=73;
sine[13095]=73;
sine[13096]=73;
sine[13097]=73;
sine[13098]=73;
sine[13099]=73;
sine[13100]=73;
sine[13101]=73;
sine[13102]=73;
sine[13103]=73;
sine[13104]=73;
sine[13105]=73;
sine[13106]=73;
sine[13107]=73;
sine[13108]=72;
sine[13109]=72;
sine[13110]=72;
sine[13111]=72;
sine[13112]=72;
sine[13113]=72;
sine[13114]=72;
sine[13115]=72;
sine[13116]=72;
sine[13117]=72;
sine[13118]=72;
sine[13119]=72;
sine[13120]=72;
sine[13121]=72;
sine[13122]=72;
sine[13123]=72;
sine[13124]=72;
sine[13125]=72;
sine[13126]=72;
sine[13127]=72;
sine[13128]=72;
sine[13129]=72;
sine[13130]=72;
sine[13131]=72;
sine[13132]=72;
sine[13133]=72;
sine[13134]=72;
sine[13135]=72;
sine[13136]=72;
sine[13137]=72;
sine[13138]=72;
sine[13139]=72;
sine[13140]=72;
sine[13141]=72;
sine[13142]=72;
sine[13143]=72;
sine[13144]=72;
sine[13145]=72;
sine[13146]=72;
sine[13147]=72;
sine[13148]=72;
sine[13149]=72;
sine[13150]=72;
sine[13151]=72;
sine[13152]=72;
sine[13153]=72;
sine[13154]=72;
sine[13155]=72;
sine[13156]=72;
sine[13157]=72;
sine[13158]=72;
sine[13159]=72;
sine[13160]=72;
sine[13161]=71;
sine[13162]=71;
sine[13163]=71;
sine[13164]=71;
sine[13165]=71;
sine[13166]=71;
sine[13167]=71;
sine[13168]=71;
sine[13169]=71;
sine[13170]=71;
sine[13171]=71;
sine[13172]=71;
sine[13173]=71;
sine[13174]=71;
sine[13175]=71;
sine[13176]=71;
sine[13177]=71;
sine[13178]=71;
sine[13179]=71;
sine[13180]=71;
sine[13181]=71;
sine[13182]=71;
sine[13183]=71;
sine[13184]=71;
sine[13185]=71;
sine[13186]=71;
sine[13187]=71;
sine[13188]=71;
sine[13189]=71;
sine[13190]=71;
sine[13191]=71;
sine[13192]=71;
sine[13193]=71;
sine[13194]=71;
sine[13195]=71;
sine[13196]=71;
sine[13197]=71;
sine[13198]=71;
sine[13199]=71;
sine[13200]=71;
sine[13201]=71;
sine[13202]=71;
sine[13203]=71;
sine[13204]=71;
sine[13205]=71;
sine[13206]=71;
sine[13207]=71;
sine[13208]=71;
sine[13209]=71;
sine[13210]=70;
sine[13211]=70;
sine[13212]=70;
sine[13213]=70;
sine[13214]=70;
sine[13215]=70;
sine[13216]=70;
sine[13217]=70;
sine[13218]=70;
sine[13219]=70;
sine[13220]=70;
sine[13221]=70;
sine[13222]=70;
sine[13223]=70;
sine[13224]=70;
sine[13225]=70;
sine[13226]=70;
sine[13227]=70;
sine[13228]=70;
sine[13229]=70;
sine[13230]=70;
sine[13231]=70;
sine[13232]=70;
sine[13233]=70;
sine[13234]=70;
sine[13235]=70;
sine[13236]=70;
sine[13237]=70;
sine[13238]=70;
sine[13239]=70;
sine[13240]=70;
sine[13241]=70;
sine[13242]=70;
sine[13243]=70;
sine[13244]=70;
sine[13245]=70;
sine[13246]=70;
sine[13247]=70;
sine[13248]=70;
sine[13249]=70;
sine[13250]=70;
sine[13251]=70;
sine[13252]=70;
sine[13253]=70;
sine[13254]=70;
sine[13255]=69;
sine[13256]=69;
sine[13257]=69;
sine[13258]=69;
sine[13259]=69;
sine[13260]=69;
sine[13261]=69;
sine[13262]=69;
sine[13263]=69;
sine[13264]=69;
sine[13265]=69;
sine[13266]=69;
sine[13267]=69;
sine[13268]=69;
sine[13269]=69;
sine[13270]=69;
sine[13271]=69;
sine[13272]=69;
sine[13273]=69;
sine[13274]=69;
sine[13275]=69;
sine[13276]=69;
sine[13277]=69;
sine[13278]=69;
sine[13279]=69;
sine[13280]=69;
sine[13281]=69;
sine[13282]=69;
sine[13283]=69;
sine[13284]=69;
sine[13285]=69;
sine[13286]=69;
sine[13287]=69;
sine[13288]=69;
sine[13289]=69;
sine[13290]=69;
sine[13291]=69;
sine[13292]=69;
sine[13293]=69;
sine[13294]=69;
sine[13295]=69;
sine[13296]=69;
sine[13297]=69;
sine[13298]=69;
sine[13299]=68;
sine[13300]=68;
sine[13301]=68;
sine[13302]=68;
sine[13303]=68;
sine[13304]=68;
sine[13305]=68;
sine[13306]=68;
sine[13307]=68;
sine[13308]=68;
sine[13309]=68;
sine[13310]=68;
sine[13311]=68;
sine[13312]=68;
sine[13313]=68;
sine[13314]=68;
sine[13315]=68;
sine[13316]=68;
sine[13317]=68;
sine[13318]=68;
sine[13319]=68;
sine[13320]=68;
sine[13321]=68;
sine[13322]=68;
sine[13323]=68;
sine[13324]=68;
sine[13325]=68;
sine[13326]=68;
sine[13327]=68;
sine[13328]=68;
sine[13329]=68;
sine[13330]=68;
sine[13331]=68;
sine[13332]=68;
sine[13333]=68;
sine[13334]=68;
sine[13335]=68;
sine[13336]=68;
sine[13337]=68;
sine[13338]=68;
sine[13339]=68;
sine[13340]=67;
sine[13341]=67;
sine[13342]=67;
sine[13343]=67;
sine[13344]=67;
sine[13345]=67;
sine[13346]=67;
sine[13347]=67;
sine[13348]=67;
sine[13349]=67;
sine[13350]=67;
sine[13351]=67;
sine[13352]=67;
sine[13353]=67;
sine[13354]=67;
sine[13355]=67;
sine[13356]=67;
sine[13357]=67;
sine[13358]=67;
sine[13359]=67;
sine[13360]=67;
sine[13361]=67;
sine[13362]=67;
sine[13363]=67;
sine[13364]=67;
sine[13365]=67;
sine[13366]=67;
sine[13367]=67;
sine[13368]=67;
sine[13369]=67;
sine[13370]=67;
sine[13371]=67;
sine[13372]=67;
sine[13373]=67;
sine[13374]=67;
sine[13375]=67;
sine[13376]=67;
sine[13377]=67;
sine[13378]=67;
sine[13379]=67;
sine[13380]=66;
sine[13381]=66;
sine[13382]=66;
sine[13383]=66;
sine[13384]=66;
sine[13385]=66;
sine[13386]=66;
sine[13387]=66;
sine[13388]=66;
sine[13389]=66;
sine[13390]=66;
sine[13391]=66;
sine[13392]=66;
sine[13393]=66;
sine[13394]=66;
sine[13395]=66;
sine[13396]=66;
sine[13397]=66;
sine[13398]=66;
sine[13399]=66;
sine[13400]=66;
sine[13401]=66;
sine[13402]=66;
sine[13403]=66;
sine[13404]=66;
sine[13405]=66;
sine[13406]=66;
sine[13407]=66;
sine[13408]=66;
sine[13409]=66;
sine[13410]=66;
sine[13411]=66;
sine[13412]=66;
sine[13413]=66;
sine[13414]=66;
sine[13415]=66;
sine[13416]=66;
sine[13417]=66;
sine[13418]=65;
sine[13419]=65;
sine[13420]=65;
sine[13421]=65;
sine[13422]=65;
sine[13423]=65;
sine[13424]=65;
sine[13425]=65;
sine[13426]=65;
sine[13427]=65;
sine[13428]=65;
sine[13429]=65;
sine[13430]=65;
sine[13431]=65;
sine[13432]=65;
sine[13433]=65;
sine[13434]=65;
sine[13435]=65;
sine[13436]=65;
sine[13437]=65;
sine[13438]=65;
sine[13439]=65;
sine[13440]=65;
sine[13441]=65;
sine[13442]=65;
sine[13443]=65;
sine[13444]=65;
sine[13445]=65;
sine[13446]=65;
sine[13447]=65;
sine[13448]=65;
sine[13449]=65;
sine[13450]=65;
sine[13451]=65;
sine[13452]=65;
sine[13453]=65;
sine[13454]=65;
sine[13455]=64;
sine[13456]=64;
sine[13457]=64;
sine[13458]=64;
sine[13459]=64;
sine[13460]=64;
sine[13461]=64;
sine[13462]=64;
sine[13463]=64;
sine[13464]=64;
sine[13465]=64;
sine[13466]=64;
sine[13467]=64;
sine[13468]=64;
sine[13469]=64;
sine[13470]=64;
sine[13471]=64;
sine[13472]=64;
sine[13473]=64;
sine[13474]=64;
sine[13475]=64;
sine[13476]=64;
sine[13477]=64;
sine[13478]=64;
sine[13479]=64;
sine[13480]=64;
sine[13481]=64;
sine[13482]=64;
sine[13483]=64;
sine[13484]=64;
sine[13485]=64;
sine[13486]=64;
sine[13487]=64;
sine[13488]=64;
sine[13489]=64;
sine[13490]=63;
sine[13491]=63;
sine[13492]=63;
sine[13493]=63;
sine[13494]=63;
sine[13495]=63;
sine[13496]=63;
sine[13497]=63;
sine[13498]=63;
sine[13499]=63;
sine[13500]=63;
sine[13501]=63;
sine[13502]=63;
sine[13503]=63;
sine[13504]=63;
sine[13505]=63;
sine[13506]=63;
sine[13507]=63;
sine[13508]=63;
sine[13509]=63;
sine[13510]=63;
sine[13511]=63;
sine[13512]=63;
sine[13513]=63;
sine[13514]=63;
sine[13515]=63;
sine[13516]=63;
sine[13517]=63;
sine[13518]=63;
sine[13519]=63;
sine[13520]=63;
sine[13521]=63;
sine[13522]=63;
sine[13523]=63;
sine[13524]=63;
sine[13525]=62;
sine[13526]=62;
sine[13527]=62;
sine[13528]=62;
sine[13529]=62;
sine[13530]=62;
sine[13531]=62;
sine[13532]=62;
sine[13533]=62;
sine[13534]=62;
sine[13535]=62;
sine[13536]=62;
sine[13537]=62;
sine[13538]=62;
sine[13539]=62;
sine[13540]=62;
sine[13541]=62;
sine[13542]=62;
sine[13543]=62;
sine[13544]=62;
sine[13545]=62;
sine[13546]=62;
sine[13547]=62;
sine[13548]=62;
sine[13549]=62;
sine[13550]=62;
sine[13551]=62;
sine[13552]=62;
sine[13553]=62;
sine[13554]=62;
sine[13555]=62;
sine[13556]=62;
sine[13557]=62;
sine[13558]=61;
sine[13559]=61;
sine[13560]=61;
sine[13561]=61;
sine[13562]=61;
sine[13563]=61;
sine[13564]=61;
sine[13565]=61;
sine[13566]=61;
sine[13567]=61;
sine[13568]=61;
sine[13569]=61;
sine[13570]=61;
sine[13571]=61;
sine[13572]=61;
sine[13573]=61;
sine[13574]=61;
sine[13575]=61;
sine[13576]=61;
sine[13577]=61;
sine[13578]=61;
sine[13579]=61;
sine[13580]=61;
sine[13581]=61;
sine[13582]=61;
sine[13583]=61;
sine[13584]=61;
sine[13585]=61;
sine[13586]=61;
sine[13587]=61;
sine[13588]=61;
sine[13589]=61;
sine[13590]=61;
sine[13591]=60;
sine[13592]=60;
sine[13593]=60;
sine[13594]=60;
sine[13595]=60;
sine[13596]=60;
sine[13597]=60;
sine[13598]=60;
sine[13599]=60;
sine[13600]=60;
sine[13601]=60;
sine[13602]=60;
sine[13603]=60;
sine[13604]=60;
sine[13605]=60;
sine[13606]=60;
sine[13607]=60;
sine[13608]=60;
sine[13609]=60;
sine[13610]=60;
sine[13611]=60;
sine[13612]=60;
sine[13613]=60;
sine[13614]=60;
sine[13615]=60;
sine[13616]=60;
sine[13617]=60;
sine[13618]=60;
sine[13619]=60;
sine[13620]=60;
sine[13621]=60;
sine[13622]=60;
sine[13623]=59;
sine[13624]=59;
sine[13625]=59;
sine[13626]=59;
sine[13627]=59;
sine[13628]=59;
sine[13629]=59;
sine[13630]=59;
sine[13631]=59;
sine[13632]=59;
sine[13633]=59;
sine[13634]=59;
sine[13635]=59;
sine[13636]=59;
sine[13637]=59;
sine[13638]=59;
sine[13639]=59;
sine[13640]=59;
sine[13641]=59;
sine[13642]=59;
sine[13643]=59;
sine[13644]=59;
sine[13645]=59;
sine[13646]=59;
sine[13647]=59;
sine[13648]=59;
sine[13649]=59;
sine[13650]=59;
sine[13651]=59;
sine[13652]=59;
sine[13653]=59;
sine[13654]=58;
sine[13655]=58;
sine[13656]=58;
sine[13657]=58;
sine[13658]=58;
sine[13659]=58;
sine[13660]=58;
sine[13661]=58;
sine[13662]=58;
sine[13663]=58;
sine[13664]=58;
sine[13665]=58;
sine[13666]=58;
sine[13667]=58;
sine[13668]=58;
sine[13669]=58;
sine[13670]=58;
sine[13671]=58;
sine[13672]=58;
sine[13673]=58;
sine[13674]=58;
sine[13675]=58;
sine[13676]=58;
sine[13677]=58;
sine[13678]=58;
sine[13679]=58;
sine[13680]=58;
sine[13681]=58;
sine[13682]=58;
sine[13683]=58;
sine[13684]=57;
sine[13685]=57;
sine[13686]=57;
sine[13687]=57;
sine[13688]=57;
sine[13689]=57;
sine[13690]=57;
sine[13691]=57;
sine[13692]=57;
sine[13693]=57;
sine[13694]=57;
sine[13695]=57;
sine[13696]=57;
sine[13697]=57;
sine[13698]=57;
sine[13699]=57;
sine[13700]=57;
sine[13701]=57;
sine[13702]=57;
sine[13703]=57;
sine[13704]=57;
sine[13705]=57;
sine[13706]=57;
sine[13707]=57;
sine[13708]=57;
sine[13709]=57;
sine[13710]=57;
sine[13711]=57;
sine[13712]=57;
sine[13713]=57;
sine[13714]=56;
sine[13715]=56;
sine[13716]=56;
sine[13717]=56;
sine[13718]=56;
sine[13719]=56;
sine[13720]=56;
sine[13721]=56;
sine[13722]=56;
sine[13723]=56;
sine[13724]=56;
sine[13725]=56;
sine[13726]=56;
sine[13727]=56;
sine[13728]=56;
sine[13729]=56;
sine[13730]=56;
sine[13731]=56;
sine[13732]=56;
sine[13733]=56;
sine[13734]=56;
sine[13735]=56;
sine[13736]=56;
sine[13737]=56;
sine[13738]=56;
sine[13739]=56;
sine[13740]=56;
sine[13741]=56;
sine[13742]=56;
sine[13743]=55;
sine[13744]=55;
sine[13745]=55;
sine[13746]=55;
sine[13747]=55;
sine[13748]=55;
sine[13749]=55;
sine[13750]=55;
sine[13751]=55;
sine[13752]=55;
sine[13753]=55;
sine[13754]=55;
sine[13755]=55;
sine[13756]=55;
sine[13757]=55;
sine[13758]=55;
sine[13759]=55;
sine[13760]=55;
sine[13761]=55;
sine[13762]=55;
sine[13763]=55;
sine[13764]=55;
sine[13765]=55;
sine[13766]=55;
sine[13767]=55;
sine[13768]=55;
sine[13769]=55;
sine[13770]=55;
sine[13771]=55;
sine[13772]=54;
sine[13773]=54;
sine[13774]=54;
sine[13775]=54;
sine[13776]=54;
sine[13777]=54;
sine[13778]=54;
sine[13779]=54;
sine[13780]=54;
sine[13781]=54;
sine[13782]=54;
sine[13783]=54;
sine[13784]=54;
sine[13785]=54;
sine[13786]=54;
sine[13787]=54;
sine[13788]=54;
sine[13789]=54;
sine[13790]=54;
sine[13791]=54;
sine[13792]=54;
sine[13793]=54;
sine[13794]=54;
sine[13795]=54;
sine[13796]=54;
sine[13797]=54;
sine[13798]=54;
sine[13799]=54;
sine[13800]=53;
sine[13801]=53;
sine[13802]=53;
sine[13803]=53;
sine[13804]=53;
sine[13805]=53;
sine[13806]=53;
sine[13807]=53;
sine[13808]=53;
sine[13809]=53;
sine[13810]=53;
sine[13811]=53;
sine[13812]=53;
sine[13813]=53;
sine[13814]=53;
sine[13815]=53;
sine[13816]=53;
sine[13817]=53;
sine[13818]=53;
sine[13819]=53;
sine[13820]=53;
sine[13821]=53;
sine[13822]=53;
sine[13823]=53;
sine[13824]=53;
sine[13825]=53;
sine[13826]=53;
sine[13827]=53;
sine[13828]=52;
sine[13829]=52;
sine[13830]=52;
sine[13831]=52;
sine[13832]=52;
sine[13833]=52;
sine[13834]=52;
sine[13835]=52;
sine[13836]=52;
sine[13837]=52;
sine[13838]=52;
sine[13839]=52;
sine[13840]=52;
sine[13841]=52;
sine[13842]=52;
sine[13843]=52;
sine[13844]=52;
sine[13845]=52;
sine[13846]=52;
sine[13847]=52;
sine[13848]=52;
sine[13849]=52;
sine[13850]=52;
sine[13851]=52;
sine[13852]=52;
sine[13853]=52;
sine[13854]=52;
sine[13855]=51;
sine[13856]=51;
sine[13857]=51;
sine[13858]=51;
sine[13859]=51;
sine[13860]=51;
sine[13861]=51;
sine[13862]=51;
sine[13863]=51;
sine[13864]=51;
sine[13865]=51;
sine[13866]=51;
sine[13867]=51;
sine[13868]=51;
sine[13869]=51;
sine[13870]=51;
sine[13871]=51;
sine[13872]=51;
sine[13873]=51;
sine[13874]=51;
sine[13875]=51;
sine[13876]=51;
sine[13877]=51;
sine[13878]=51;
sine[13879]=51;
sine[13880]=51;
sine[13881]=51;
sine[13882]=50;
sine[13883]=50;
sine[13884]=50;
sine[13885]=50;
sine[13886]=50;
sine[13887]=50;
sine[13888]=50;
sine[13889]=50;
sine[13890]=50;
sine[13891]=50;
sine[13892]=50;
sine[13893]=50;
sine[13894]=50;
sine[13895]=50;
sine[13896]=50;
sine[13897]=50;
sine[13898]=50;
sine[13899]=50;
sine[13900]=50;
sine[13901]=50;
sine[13902]=50;
sine[13903]=50;
sine[13904]=50;
sine[13905]=50;
sine[13906]=50;
sine[13907]=50;
sine[13908]=49;
sine[13909]=49;
sine[13910]=49;
sine[13911]=49;
sine[13912]=49;
sine[13913]=49;
sine[13914]=49;
sine[13915]=49;
sine[13916]=49;
sine[13917]=49;
sine[13918]=49;
sine[13919]=49;
sine[13920]=49;
sine[13921]=49;
sine[13922]=49;
sine[13923]=49;
sine[13924]=49;
sine[13925]=49;
sine[13926]=49;
sine[13927]=49;
sine[13928]=49;
sine[13929]=49;
sine[13930]=49;
sine[13931]=49;
sine[13932]=49;
sine[13933]=49;
sine[13934]=49;
sine[13935]=48;
sine[13936]=48;
sine[13937]=48;
sine[13938]=48;
sine[13939]=48;
sine[13940]=48;
sine[13941]=48;
sine[13942]=48;
sine[13943]=48;
sine[13944]=48;
sine[13945]=48;
sine[13946]=48;
sine[13947]=48;
sine[13948]=48;
sine[13949]=48;
sine[13950]=48;
sine[13951]=48;
sine[13952]=48;
sine[13953]=48;
sine[13954]=48;
sine[13955]=48;
sine[13956]=48;
sine[13957]=48;
sine[13958]=48;
sine[13959]=48;
sine[13960]=47;
sine[13961]=47;
sine[13962]=47;
sine[13963]=47;
sine[13964]=47;
sine[13965]=47;
sine[13966]=47;
sine[13967]=47;
sine[13968]=47;
sine[13969]=47;
sine[13970]=47;
sine[13971]=47;
sine[13972]=47;
sine[13973]=47;
sine[13974]=47;
sine[13975]=47;
sine[13976]=47;
sine[13977]=47;
sine[13978]=47;
sine[13979]=47;
sine[13980]=47;
sine[13981]=47;
sine[13982]=47;
sine[13983]=47;
sine[13984]=47;
sine[13985]=47;
sine[13986]=46;
sine[13987]=46;
sine[13988]=46;
sine[13989]=46;
sine[13990]=46;
sine[13991]=46;
sine[13992]=46;
sine[13993]=46;
sine[13994]=46;
sine[13995]=46;
sine[13996]=46;
sine[13997]=46;
sine[13998]=46;
sine[13999]=46;
sine[14000]=46;
sine[14001]=46;
sine[14002]=46;
sine[14003]=46;
sine[14004]=46;
sine[14005]=46;
sine[14006]=46;
sine[14007]=46;
sine[14008]=46;
sine[14009]=46;
sine[14010]=46;
sine[14011]=45;
sine[14012]=45;
sine[14013]=45;
sine[14014]=45;
sine[14015]=45;
sine[14016]=45;
sine[14017]=45;
sine[14018]=45;
sine[14019]=45;
sine[14020]=45;
sine[14021]=45;
sine[14022]=45;
sine[14023]=45;
sine[14024]=45;
sine[14025]=45;
sine[14026]=45;
sine[14027]=45;
sine[14028]=45;
sine[14029]=45;
sine[14030]=45;
sine[14031]=45;
sine[14032]=45;
sine[14033]=45;
sine[14034]=45;
sine[14035]=45;
sine[14036]=44;
sine[14037]=44;
sine[14038]=44;
sine[14039]=44;
sine[14040]=44;
sine[14041]=44;
sine[14042]=44;
sine[14043]=44;
sine[14044]=44;
sine[14045]=44;
sine[14046]=44;
sine[14047]=44;
sine[14048]=44;
sine[14049]=44;
sine[14050]=44;
sine[14051]=44;
sine[14052]=44;
sine[14053]=44;
sine[14054]=44;
sine[14055]=44;
sine[14056]=44;
sine[14057]=44;
sine[14058]=44;
sine[14059]=44;
sine[14060]=44;
sine[14061]=43;
sine[14062]=43;
sine[14063]=43;
sine[14064]=43;
sine[14065]=43;
sine[14066]=43;
sine[14067]=43;
sine[14068]=43;
sine[14069]=43;
sine[14070]=43;
sine[14071]=43;
sine[14072]=43;
sine[14073]=43;
sine[14074]=43;
sine[14075]=43;
sine[14076]=43;
sine[14077]=43;
sine[14078]=43;
sine[14079]=43;
sine[14080]=43;
sine[14081]=43;
sine[14082]=43;
sine[14083]=43;
sine[14084]=43;
sine[14085]=42;
sine[14086]=42;
sine[14087]=42;
sine[14088]=42;
sine[14089]=42;
sine[14090]=42;
sine[14091]=42;
sine[14092]=42;
sine[14093]=42;
sine[14094]=42;
sine[14095]=42;
sine[14096]=42;
sine[14097]=42;
sine[14098]=42;
sine[14099]=42;
sine[14100]=42;
sine[14101]=42;
sine[14102]=42;
sine[14103]=42;
sine[14104]=42;
sine[14105]=42;
sine[14106]=42;
sine[14107]=42;
sine[14108]=42;
sine[14109]=41;
sine[14110]=41;
sine[14111]=41;
sine[14112]=41;
sine[14113]=41;
sine[14114]=41;
sine[14115]=41;
sine[14116]=41;
sine[14117]=41;
sine[14118]=41;
sine[14119]=41;
sine[14120]=41;
sine[14121]=41;
sine[14122]=41;
sine[14123]=41;
sine[14124]=41;
sine[14125]=41;
sine[14126]=41;
sine[14127]=41;
sine[14128]=41;
sine[14129]=41;
sine[14130]=41;
sine[14131]=41;
sine[14132]=41;
sine[14133]=40;
sine[14134]=40;
sine[14135]=40;
sine[14136]=40;
sine[14137]=40;
sine[14138]=40;
sine[14139]=40;
sine[14140]=40;
sine[14141]=40;
sine[14142]=40;
sine[14143]=40;
sine[14144]=40;
sine[14145]=40;
sine[14146]=40;
sine[14147]=40;
sine[14148]=40;
sine[14149]=40;
sine[14150]=40;
sine[14151]=40;
sine[14152]=40;
sine[14153]=40;
sine[14154]=40;
sine[14155]=40;
sine[14156]=40;
sine[14157]=39;
sine[14158]=39;
sine[14159]=39;
sine[14160]=39;
sine[14161]=39;
sine[14162]=39;
sine[14163]=39;
sine[14164]=39;
sine[14165]=39;
sine[14166]=39;
sine[14167]=39;
sine[14168]=39;
sine[14169]=39;
sine[14170]=39;
sine[14171]=39;
sine[14172]=39;
sine[14173]=39;
sine[14174]=39;
sine[14175]=39;
sine[14176]=39;
sine[14177]=39;
sine[14178]=39;
sine[14179]=39;
sine[14180]=38;
sine[14181]=38;
sine[14182]=38;
sine[14183]=38;
sine[14184]=38;
sine[14185]=38;
sine[14186]=38;
sine[14187]=38;
sine[14188]=38;
sine[14189]=38;
sine[14190]=38;
sine[14191]=38;
sine[14192]=38;
sine[14193]=38;
sine[14194]=38;
sine[14195]=38;
sine[14196]=38;
sine[14197]=38;
sine[14198]=38;
sine[14199]=38;
sine[14200]=38;
sine[14201]=38;
sine[14202]=38;
sine[14203]=38;
sine[14204]=37;
sine[14205]=37;
sine[14206]=37;
sine[14207]=37;
sine[14208]=37;
sine[14209]=37;
sine[14210]=37;
sine[14211]=37;
sine[14212]=37;
sine[14213]=37;
sine[14214]=37;
sine[14215]=37;
sine[14216]=37;
sine[14217]=37;
sine[14218]=37;
sine[14219]=37;
sine[14220]=37;
sine[14221]=37;
sine[14222]=37;
sine[14223]=37;
sine[14224]=37;
sine[14225]=37;
sine[14226]=37;
sine[14227]=36;
sine[14228]=36;
sine[14229]=36;
sine[14230]=36;
sine[14231]=36;
sine[14232]=36;
sine[14233]=36;
sine[14234]=36;
sine[14235]=36;
sine[14236]=36;
sine[14237]=36;
sine[14238]=36;
sine[14239]=36;
sine[14240]=36;
sine[14241]=36;
sine[14242]=36;
sine[14243]=36;
sine[14244]=36;
sine[14245]=36;
sine[14246]=36;
sine[14247]=36;
sine[14248]=36;
sine[14249]=36;
sine[14250]=35;
sine[14251]=35;
sine[14252]=35;
sine[14253]=35;
sine[14254]=35;
sine[14255]=35;
sine[14256]=35;
sine[14257]=35;
sine[14258]=35;
sine[14259]=35;
sine[14260]=35;
sine[14261]=35;
sine[14262]=35;
sine[14263]=35;
sine[14264]=35;
sine[14265]=35;
sine[14266]=35;
sine[14267]=35;
sine[14268]=35;
sine[14269]=35;
sine[14270]=35;
sine[14271]=35;
sine[14272]=35;
sine[14273]=34;
sine[14274]=34;
sine[14275]=34;
sine[14276]=34;
sine[14277]=34;
sine[14278]=34;
sine[14279]=34;
sine[14280]=34;
sine[14281]=34;
sine[14282]=34;
sine[14283]=34;
sine[14284]=34;
sine[14285]=34;
sine[14286]=34;
sine[14287]=34;
sine[14288]=34;
sine[14289]=34;
sine[14290]=34;
sine[14291]=34;
sine[14292]=34;
sine[14293]=34;
sine[14294]=34;
sine[14295]=33;
sine[14296]=33;
sine[14297]=33;
sine[14298]=33;
sine[14299]=33;
sine[14300]=33;
sine[14301]=33;
sine[14302]=33;
sine[14303]=33;
sine[14304]=33;
sine[14305]=33;
sine[14306]=33;
sine[14307]=33;
sine[14308]=33;
sine[14309]=33;
sine[14310]=33;
sine[14311]=33;
sine[14312]=33;
sine[14313]=33;
sine[14314]=33;
sine[14315]=33;
sine[14316]=33;
sine[14317]=33;
sine[14318]=32;
sine[14319]=32;
sine[14320]=32;
sine[14321]=32;
sine[14322]=32;
sine[14323]=32;
sine[14324]=32;
sine[14325]=32;
sine[14326]=32;
sine[14327]=32;
sine[14328]=32;
sine[14329]=32;
sine[14330]=32;
sine[14331]=32;
sine[14332]=32;
sine[14333]=32;
sine[14334]=32;
sine[14335]=32;
sine[14336]=32;
sine[14337]=32;
sine[14338]=32;
sine[14339]=32;
sine[14340]=31;
sine[14341]=31;
sine[14342]=31;
sine[14343]=31;
sine[14344]=31;
sine[14345]=31;
sine[14346]=31;
sine[14347]=31;
sine[14348]=31;
sine[14349]=31;
sine[14350]=31;
sine[14351]=31;
sine[14352]=31;
sine[14353]=31;
sine[14354]=31;
sine[14355]=31;
sine[14356]=31;
sine[14357]=31;
sine[14358]=31;
sine[14359]=31;
sine[14360]=31;
sine[14361]=31;
sine[14362]=30;
sine[14363]=30;
sine[14364]=30;
sine[14365]=30;
sine[14366]=30;
sine[14367]=30;
sine[14368]=30;
sine[14369]=30;
sine[14370]=30;
sine[14371]=30;
sine[14372]=30;
sine[14373]=30;
sine[14374]=30;
sine[14375]=30;
sine[14376]=30;
sine[14377]=30;
sine[14378]=30;
sine[14379]=30;
sine[14380]=30;
sine[14381]=30;
sine[14382]=30;
sine[14383]=30;
sine[14384]=29;
sine[14385]=29;
sine[14386]=29;
sine[14387]=29;
sine[14388]=29;
sine[14389]=29;
sine[14390]=29;
sine[14391]=29;
sine[14392]=29;
sine[14393]=29;
sine[14394]=29;
sine[14395]=29;
sine[14396]=29;
sine[14397]=29;
sine[14398]=29;
sine[14399]=29;
sine[14400]=29;
sine[14401]=29;
sine[14402]=29;
sine[14403]=29;
sine[14404]=29;
sine[14405]=29;
sine[14406]=28;
sine[14407]=28;
sine[14408]=28;
sine[14409]=28;
sine[14410]=28;
sine[14411]=28;
sine[14412]=28;
sine[14413]=28;
sine[14414]=28;
sine[14415]=28;
sine[14416]=28;
sine[14417]=28;
sine[14418]=28;
sine[14419]=28;
sine[14420]=28;
sine[14421]=28;
sine[14422]=28;
sine[14423]=28;
sine[14424]=28;
sine[14425]=28;
sine[14426]=28;
sine[14427]=28;
sine[14428]=27;
sine[14429]=27;
sine[14430]=27;
sine[14431]=27;
sine[14432]=27;
sine[14433]=27;
sine[14434]=27;
sine[14435]=27;
sine[14436]=27;
sine[14437]=27;
sine[14438]=27;
sine[14439]=27;
sine[14440]=27;
sine[14441]=27;
sine[14442]=27;
sine[14443]=27;
sine[14444]=27;
sine[14445]=27;
sine[14446]=27;
sine[14447]=27;
sine[14448]=27;
sine[14449]=27;
sine[14450]=26;
sine[14451]=26;
sine[14452]=26;
sine[14453]=26;
sine[14454]=26;
sine[14455]=26;
sine[14456]=26;
sine[14457]=26;
sine[14458]=26;
sine[14459]=26;
sine[14460]=26;
sine[14461]=26;
sine[14462]=26;
sine[14463]=26;
sine[14464]=26;
sine[14465]=26;
sine[14466]=26;
sine[14467]=26;
sine[14468]=26;
sine[14469]=26;
sine[14470]=26;
sine[14471]=25;
sine[14472]=25;
sine[14473]=25;
sine[14474]=25;
sine[14475]=25;
sine[14476]=25;
sine[14477]=25;
sine[14478]=25;
sine[14479]=25;
sine[14480]=25;
sine[14481]=25;
sine[14482]=25;
sine[14483]=25;
sine[14484]=25;
sine[14485]=25;
sine[14486]=25;
sine[14487]=25;
sine[14488]=25;
sine[14489]=25;
sine[14490]=25;
sine[14491]=25;
sine[14492]=25;
sine[14493]=24;
sine[14494]=24;
sine[14495]=24;
sine[14496]=24;
sine[14497]=24;
sine[14498]=24;
sine[14499]=24;
sine[14500]=24;
sine[14501]=24;
sine[14502]=24;
sine[14503]=24;
sine[14504]=24;
sine[14505]=24;
sine[14506]=24;
sine[14507]=24;
sine[14508]=24;
sine[14509]=24;
sine[14510]=24;
sine[14511]=24;
sine[14512]=24;
sine[14513]=24;
sine[14514]=23;
sine[14515]=23;
sine[14516]=23;
sine[14517]=23;
sine[14518]=23;
sine[14519]=23;
sine[14520]=23;
sine[14521]=23;
sine[14522]=23;
sine[14523]=23;
sine[14524]=23;
sine[14525]=23;
sine[14526]=23;
sine[14527]=23;
sine[14528]=23;
sine[14529]=23;
sine[14530]=23;
sine[14531]=23;
sine[14532]=23;
sine[14533]=23;
sine[14534]=23;
sine[14535]=23;
sine[14536]=22;
sine[14537]=22;
sine[14538]=22;
sine[14539]=22;
sine[14540]=22;
sine[14541]=22;
sine[14542]=22;
sine[14543]=22;
sine[14544]=22;
sine[14545]=22;
sine[14546]=22;
sine[14547]=22;
sine[14548]=22;
sine[14549]=22;
sine[14550]=22;
sine[14551]=22;
sine[14552]=22;
sine[14553]=22;
sine[14554]=22;
sine[14555]=22;
sine[14556]=22;
sine[14557]=21;
sine[14558]=21;
sine[14559]=21;
sine[14560]=21;
sine[14561]=21;
sine[14562]=21;
sine[14563]=21;
sine[14564]=21;
sine[14565]=21;
sine[14566]=21;
sine[14567]=21;
sine[14568]=21;
sine[14569]=21;
sine[14570]=21;
sine[14571]=21;
sine[14572]=21;
sine[14573]=21;
sine[14574]=21;
sine[14575]=21;
sine[14576]=21;
sine[14577]=21;
sine[14578]=20;
sine[14579]=20;
sine[14580]=20;
sine[14581]=20;
sine[14582]=20;
sine[14583]=20;
sine[14584]=20;
sine[14585]=20;
sine[14586]=20;
sine[14587]=20;
sine[14588]=20;
sine[14589]=20;
sine[14590]=20;
sine[14591]=20;
sine[14592]=20;
sine[14593]=20;
sine[14594]=20;
sine[14595]=20;
sine[14596]=20;
sine[14597]=20;
sine[14598]=20;
sine[14599]=19;
sine[14600]=19;
sine[14601]=19;
sine[14602]=19;
sine[14603]=19;
sine[14604]=19;
sine[14605]=19;
sine[14606]=19;
sine[14607]=19;
sine[14608]=19;
sine[14609]=19;
sine[14610]=19;
sine[14611]=19;
sine[14612]=19;
sine[14613]=19;
sine[14614]=19;
sine[14615]=19;
sine[14616]=19;
sine[14617]=19;
sine[14618]=19;
sine[14619]=19;
sine[14620]=18;
sine[14621]=18;
sine[14622]=18;
sine[14623]=18;
sine[14624]=18;
sine[14625]=18;
sine[14626]=18;
sine[14627]=18;
sine[14628]=18;
sine[14629]=18;
sine[14630]=18;
sine[14631]=18;
sine[14632]=18;
sine[14633]=18;
sine[14634]=18;
sine[14635]=18;
sine[14636]=18;
sine[14637]=18;
sine[14638]=18;
sine[14639]=18;
sine[14640]=18;
sine[14641]=17;
sine[14642]=17;
sine[14643]=17;
sine[14644]=17;
sine[14645]=17;
sine[14646]=17;
sine[14647]=17;
sine[14648]=17;
sine[14649]=17;
sine[14650]=17;
sine[14651]=17;
sine[14652]=17;
sine[14653]=17;
sine[14654]=17;
sine[14655]=17;
sine[14656]=17;
sine[14657]=17;
sine[14658]=17;
sine[14659]=17;
sine[14660]=17;
sine[14661]=17;
sine[14662]=16;
sine[14663]=16;
sine[14664]=16;
sine[14665]=16;
sine[14666]=16;
sine[14667]=16;
sine[14668]=16;
sine[14669]=16;
sine[14670]=16;
sine[14671]=16;
sine[14672]=16;
sine[14673]=16;
sine[14674]=16;
sine[14675]=16;
sine[14676]=16;
sine[14677]=16;
sine[14678]=16;
sine[14679]=16;
sine[14680]=16;
sine[14681]=16;
sine[14682]=16;
sine[14683]=15;
sine[14684]=15;
sine[14685]=15;
sine[14686]=15;
sine[14687]=15;
sine[14688]=15;
sine[14689]=15;
sine[14690]=15;
sine[14691]=15;
sine[14692]=15;
sine[14693]=15;
sine[14694]=15;
sine[14695]=15;
sine[14696]=15;
sine[14697]=15;
sine[14698]=15;
sine[14699]=15;
sine[14700]=15;
sine[14701]=15;
sine[14702]=15;
sine[14703]=14;
sine[14704]=14;
sine[14705]=14;
sine[14706]=14;
sine[14707]=14;
sine[14708]=14;
sine[14709]=14;
sine[14710]=14;
sine[14711]=14;
sine[14712]=14;
sine[14713]=14;
sine[14714]=14;
sine[14715]=14;
sine[14716]=14;
sine[14717]=14;
sine[14718]=14;
sine[14719]=14;
sine[14720]=14;
sine[14721]=14;
sine[14722]=14;
sine[14723]=14;
sine[14724]=13;
sine[14725]=13;
sine[14726]=13;
sine[14727]=13;
sine[14728]=13;
sine[14729]=13;
sine[14730]=13;
sine[14731]=13;
sine[14732]=13;
sine[14733]=13;
sine[14734]=13;
sine[14735]=13;
sine[14736]=13;
sine[14737]=13;
sine[14738]=13;
sine[14739]=13;
sine[14740]=13;
sine[14741]=13;
sine[14742]=13;
sine[14743]=13;
sine[14744]=13;
sine[14745]=12;
sine[14746]=12;
sine[14747]=12;
sine[14748]=12;
sine[14749]=12;
sine[14750]=12;
sine[14751]=12;
sine[14752]=12;
sine[14753]=12;
sine[14754]=12;
sine[14755]=12;
sine[14756]=12;
sine[14757]=12;
sine[14758]=12;
sine[14759]=12;
sine[14760]=12;
sine[14761]=12;
sine[14762]=12;
sine[14763]=12;
sine[14764]=12;
sine[14765]=11;
sine[14766]=11;
sine[14767]=11;
sine[14768]=11;
sine[14769]=11;
sine[14770]=11;
sine[14771]=11;
sine[14772]=11;
sine[14773]=11;
sine[14774]=11;
sine[14775]=11;
sine[14776]=11;
sine[14777]=11;
sine[14778]=11;
sine[14779]=11;
sine[14780]=11;
sine[14781]=11;
sine[14782]=11;
sine[14783]=11;
sine[14784]=11;
sine[14785]=11;
sine[14786]=10;
sine[14787]=10;
sine[14788]=10;
sine[14789]=10;
sine[14790]=10;
sine[14791]=10;
sine[14792]=10;
sine[14793]=10;
sine[14794]=10;
sine[14795]=10;
sine[14796]=10;
sine[14797]=10;
sine[14798]=10;
sine[14799]=10;
sine[14800]=10;
sine[14801]=10;
sine[14802]=10;
sine[14803]=10;
sine[14804]=10;
sine[14805]=10;
sine[14806]=9;
sine[14807]=9;
sine[14808]=9;
sine[14809]=9;
sine[14810]=9;
sine[14811]=9;
sine[14812]=9;
sine[14813]=9;
sine[14814]=9;
sine[14815]=9;
sine[14816]=9;
sine[14817]=9;
sine[14818]=9;
sine[14819]=9;
sine[14820]=9;
sine[14821]=9;
sine[14822]=9;
sine[14823]=9;
sine[14824]=9;
sine[14825]=9;
sine[14826]=9;
sine[14827]=8;
sine[14828]=8;
sine[14829]=8;
sine[14830]=8;
sine[14831]=8;
sine[14832]=8;
sine[14833]=8;
sine[14834]=8;
sine[14835]=8;
sine[14836]=8;
sine[14837]=8;
sine[14838]=8;
sine[14839]=8;
sine[14840]=8;
sine[14841]=8;
sine[14842]=8;
sine[14843]=8;
sine[14844]=8;
sine[14845]=8;
sine[14846]=8;
sine[14847]=7;
sine[14848]=7;
sine[14849]=7;
sine[14850]=7;
sine[14851]=7;
sine[14852]=7;
sine[14853]=7;
sine[14854]=7;
sine[14855]=7;
sine[14856]=7;
sine[14857]=7;
sine[14858]=7;
sine[14859]=7;
sine[14860]=7;
sine[14861]=7;
sine[14862]=7;
sine[14863]=7;
sine[14864]=7;
sine[14865]=7;
sine[14866]=7;
sine[14867]=7;
sine[14868]=6;
sine[14869]=6;
sine[14870]=6;
sine[14871]=6;
sine[14872]=6;
sine[14873]=6;
sine[14874]=6;
sine[14875]=6;
sine[14876]=6;
sine[14877]=6;
sine[14878]=6;
sine[14879]=6;
sine[14880]=6;
sine[14881]=6;
sine[14882]=6;
sine[14883]=6;
sine[14884]=6;
sine[14885]=6;
sine[14886]=6;
sine[14887]=6;
sine[14888]=5;
sine[14889]=5;
sine[14890]=5;
sine[14891]=5;
sine[14892]=5;
sine[14893]=5;
sine[14894]=5;
sine[14895]=5;
sine[14896]=5;
sine[14897]=5;
sine[14898]=5;
sine[14899]=5;
sine[14900]=5;
sine[14901]=5;
sine[14902]=5;
sine[14903]=5;
sine[14904]=5;
sine[14905]=5;
sine[14906]=5;
sine[14907]=5;
sine[14908]=5;
sine[14909]=4;
sine[14910]=4;
sine[14911]=4;
sine[14912]=4;
sine[14913]=4;
sine[14914]=4;
sine[14915]=4;
sine[14916]=4;
sine[14917]=4;
sine[14918]=4;
sine[14919]=4;
sine[14920]=4;
sine[14921]=4;
sine[14922]=4;
sine[14923]=4;
sine[14924]=4;
sine[14925]=4;
sine[14926]=4;
sine[14927]=4;
sine[14928]=4;
sine[14929]=3;
sine[14930]=3;
sine[14931]=3;
sine[14932]=3;
sine[14933]=3;
sine[14934]=3;
sine[14935]=3;
sine[14936]=3;
sine[14937]=3;
sine[14938]=3;
sine[14939]=3;
sine[14940]=3;
sine[14941]=3;
sine[14942]=3;
sine[14943]=3;
sine[14944]=3;
sine[14945]=3;
sine[14946]=3;
sine[14947]=3;
sine[14948]=3;
sine[14949]=3;
sine[14950]=2;
sine[14951]=2;
sine[14952]=2;
sine[14953]=2;
sine[14954]=2;
sine[14955]=2;
sine[14956]=2;
sine[14957]=2;
sine[14958]=2;
sine[14959]=2;
sine[14960]=2;
sine[14961]=2;
sine[14962]=2;
sine[14963]=2;
sine[14964]=2;
sine[14965]=2;
sine[14966]=2;
sine[14967]=2;
sine[14968]=2;
sine[14969]=2;
sine[14970]=1;
sine[14971]=1;
sine[14972]=1;
sine[14973]=1;
sine[14974]=1;
sine[14975]=1;
sine[14976]=1;
sine[14977]=1;
sine[14978]=1;
sine[14979]=1;
sine[14980]=1;
sine[14981]=1;
sine[14982]=1;
sine[14983]=1;
sine[14984]=1;
sine[14985]=1;
sine[14986]=1;
sine[14987]=1;
sine[14988]=1;
sine[14989]=1;
sine[14990]=0;
sine[14991]=0;
sine[14992]=0;
sine[14993]=0;
sine[14994]=0;
sine[14995]=0;
sine[14996]=0;
sine[14997]=0;
sine[14998]=0;
sine[14999]=0;
sine[15000]=0;
sine[15001]=0;
sine[15002]=0;
sine[15003]=0;
sine[15004]=0;
sine[15005]=0;
sine[15006]=0;
sine[15007]=0;
sine[15008]=0;
sine[15009]=0;
sine[15010]=0;
sine[15011]=-1;
sine[15012]=-1;
sine[15013]=-1;
sine[15014]=-1;
sine[15015]=-1;
sine[15016]=-1;
sine[15017]=-1;
sine[15018]=-1;
sine[15019]=-1;
sine[15020]=-1;
sine[15021]=-1;
sine[15022]=-1;
sine[15023]=-1;
sine[15024]=-1;
sine[15025]=-1;
sine[15026]=-1;
sine[15027]=-1;
sine[15028]=-1;
sine[15029]=-1;
sine[15030]=-1;
sine[15031]=-2;
sine[15032]=-2;
sine[15033]=-2;
sine[15034]=-2;
sine[15035]=-2;
sine[15036]=-2;
sine[15037]=-2;
sine[15038]=-2;
sine[15039]=-2;
sine[15040]=-2;
sine[15041]=-2;
sine[15042]=-2;
sine[15043]=-2;
sine[15044]=-2;
sine[15045]=-2;
sine[15046]=-2;
sine[15047]=-2;
sine[15048]=-2;
sine[15049]=-2;
sine[15050]=-2;
sine[15051]=-3;
sine[15052]=-3;
sine[15053]=-3;
sine[15054]=-3;
sine[15055]=-3;
sine[15056]=-3;
sine[15057]=-3;
sine[15058]=-3;
sine[15059]=-3;
sine[15060]=-3;
sine[15061]=-3;
sine[15062]=-3;
sine[15063]=-3;
sine[15064]=-3;
sine[15065]=-3;
sine[15066]=-3;
sine[15067]=-3;
sine[15068]=-3;
sine[15069]=-3;
sine[15070]=-3;
sine[15071]=-3;
sine[15072]=-4;
sine[15073]=-4;
sine[15074]=-4;
sine[15075]=-4;
sine[15076]=-4;
sine[15077]=-4;
sine[15078]=-4;
sine[15079]=-4;
sine[15080]=-4;
sine[15081]=-4;
sine[15082]=-4;
sine[15083]=-4;
sine[15084]=-4;
sine[15085]=-4;
sine[15086]=-4;
sine[15087]=-4;
sine[15088]=-4;
sine[15089]=-4;
sine[15090]=-4;
sine[15091]=-4;
sine[15092]=-5;
sine[15093]=-5;
sine[15094]=-5;
sine[15095]=-5;
sine[15096]=-5;
sine[15097]=-5;
sine[15098]=-5;
sine[15099]=-5;
sine[15100]=-5;
sine[15101]=-5;
sine[15102]=-5;
sine[15103]=-5;
sine[15104]=-5;
sine[15105]=-5;
sine[15106]=-5;
sine[15107]=-5;
sine[15108]=-5;
sine[15109]=-5;
sine[15110]=-5;
sine[15111]=-5;
sine[15112]=-5;
sine[15113]=-6;
sine[15114]=-6;
sine[15115]=-6;
sine[15116]=-6;
sine[15117]=-6;
sine[15118]=-6;
sine[15119]=-6;
sine[15120]=-6;
sine[15121]=-6;
sine[15122]=-6;
sine[15123]=-6;
sine[15124]=-6;
sine[15125]=-6;
sine[15126]=-6;
sine[15127]=-6;
sine[15128]=-6;
sine[15129]=-6;
sine[15130]=-6;
sine[15131]=-6;
sine[15132]=-6;
sine[15133]=-7;
sine[15134]=-7;
sine[15135]=-7;
sine[15136]=-7;
sine[15137]=-7;
sine[15138]=-7;
sine[15139]=-7;
sine[15140]=-7;
sine[15141]=-7;
sine[15142]=-7;
sine[15143]=-7;
sine[15144]=-7;
sine[15145]=-7;
sine[15146]=-7;
sine[15147]=-7;
sine[15148]=-7;
sine[15149]=-7;
sine[15150]=-7;
sine[15151]=-7;
sine[15152]=-7;
sine[15153]=-7;
sine[15154]=-8;
sine[15155]=-8;
sine[15156]=-8;
sine[15157]=-8;
sine[15158]=-8;
sine[15159]=-8;
sine[15160]=-8;
sine[15161]=-8;
sine[15162]=-8;
sine[15163]=-8;
sine[15164]=-8;
sine[15165]=-8;
sine[15166]=-8;
sine[15167]=-8;
sine[15168]=-8;
sine[15169]=-8;
sine[15170]=-8;
sine[15171]=-8;
sine[15172]=-8;
sine[15173]=-8;
sine[15174]=-9;
sine[15175]=-9;
sine[15176]=-9;
sine[15177]=-9;
sine[15178]=-9;
sine[15179]=-9;
sine[15180]=-9;
sine[15181]=-9;
sine[15182]=-9;
sine[15183]=-9;
sine[15184]=-9;
sine[15185]=-9;
sine[15186]=-9;
sine[15187]=-9;
sine[15188]=-9;
sine[15189]=-9;
sine[15190]=-9;
sine[15191]=-9;
sine[15192]=-9;
sine[15193]=-9;
sine[15194]=-9;
sine[15195]=-10;
sine[15196]=-10;
sine[15197]=-10;
sine[15198]=-10;
sine[15199]=-10;
sine[15200]=-10;
sine[15201]=-10;
sine[15202]=-10;
sine[15203]=-10;
sine[15204]=-10;
sine[15205]=-10;
sine[15206]=-10;
sine[15207]=-10;
sine[15208]=-10;
sine[15209]=-10;
sine[15210]=-10;
sine[15211]=-10;
sine[15212]=-10;
sine[15213]=-10;
sine[15214]=-10;
sine[15215]=-11;
sine[15216]=-11;
sine[15217]=-11;
sine[15218]=-11;
sine[15219]=-11;
sine[15220]=-11;
sine[15221]=-11;
sine[15222]=-11;
sine[15223]=-11;
sine[15224]=-11;
sine[15225]=-11;
sine[15226]=-11;
sine[15227]=-11;
sine[15228]=-11;
sine[15229]=-11;
sine[15230]=-11;
sine[15231]=-11;
sine[15232]=-11;
sine[15233]=-11;
sine[15234]=-11;
sine[15235]=-11;
sine[15236]=-12;
sine[15237]=-12;
sine[15238]=-12;
sine[15239]=-12;
sine[15240]=-12;
sine[15241]=-12;
sine[15242]=-12;
sine[15243]=-12;
sine[15244]=-12;
sine[15245]=-12;
sine[15246]=-12;
sine[15247]=-12;
sine[15248]=-12;
sine[15249]=-12;
sine[15250]=-12;
sine[15251]=-12;
sine[15252]=-12;
sine[15253]=-12;
sine[15254]=-12;
sine[15255]=-12;
sine[15256]=-13;
sine[15257]=-13;
sine[15258]=-13;
sine[15259]=-13;
sine[15260]=-13;
sine[15261]=-13;
sine[15262]=-13;
sine[15263]=-13;
sine[15264]=-13;
sine[15265]=-13;
sine[15266]=-13;
sine[15267]=-13;
sine[15268]=-13;
sine[15269]=-13;
sine[15270]=-13;
sine[15271]=-13;
sine[15272]=-13;
sine[15273]=-13;
sine[15274]=-13;
sine[15275]=-13;
sine[15276]=-13;
sine[15277]=-14;
sine[15278]=-14;
sine[15279]=-14;
sine[15280]=-14;
sine[15281]=-14;
sine[15282]=-14;
sine[15283]=-14;
sine[15284]=-14;
sine[15285]=-14;
sine[15286]=-14;
sine[15287]=-14;
sine[15288]=-14;
sine[15289]=-14;
sine[15290]=-14;
sine[15291]=-14;
sine[15292]=-14;
sine[15293]=-14;
sine[15294]=-14;
sine[15295]=-14;
sine[15296]=-14;
sine[15297]=-14;
sine[15298]=-15;
sine[15299]=-15;
sine[15300]=-15;
sine[15301]=-15;
sine[15302]=-15;
sine[15303]=-15;
sine[15304]=-15;
sine[15305]=-15;
sine[15306]=-15;
sine[15307]=-15;
sine[15308]=-15;
sine[15309]=-15;
sine[15310]=-15;
sine[15311]=-15;
sine[15312]=-15;
sine[15313]=-15;
sine[15314]=-15;
sine[15315]=-15;
sine[15316]=-15;
sine[15317]=-15;
sine[15318]=-16;
sine[15319]=-16;
sine[15320]=-16;
sine[15321]=-16;
sine[15322]=-16;
sine[15323]=-16;
sine[15324]=-16;
sine[15325]=-16;
sine[15326]=-16;
sine[15327]=-16;
sine[15328]=-16;
sine[15329]=-16;
sine[15330]=-16;
sine[15331]=-16;
sine[15332]=-16;
sine[15333]=-16;
sine[15334]=-16;
sine[15335]=-16;
sine[15336]=-16;
sine[15337]=-16;
sine[15338]=-16;
sine[15339]=-17;
sine[15340]=-17;
sine[15341]=-17;
sine[15342]=-17;
sine[15343]=-17;
sine[15344]=-17;
sine[15345]=-17;
sine[15346]=-17;
sine[15347]=-17;
sine[15348]=-17;
sine[15349]=-17;
sine[15350]=-17;
sine[15351]=-17;
sine[15352]=-17;
sine[15353]=-17;
sine[15354]=-17;
sine[15355]=-17;
sine[15356]=-17;
sine[15357]=-17;
sine[15358]=-17;
sine[15359]=-17;
sine[15360]=-18;
sine[15361]=-18;
sine[15362]=-18;
sine[15363]=-18;
sine[15364]=-18;
sine[15365]=-18;
sine[15366]=-18;
sine[15367]=-18;
sine[15368]=-18;
sine[15369]=-18;
sine[15370]=-18;
sine[15371]=-18;
sine[15372]=-18;
sine[15373]=-18;
sine[15374]=-18;
sine[15375]=-18;
sine[15376]=-18;
sine[15377]=-18;
sine[15378]=-18;
sine[15379]=-18;
sine[15380]=-18;
sine[15381]=-19;
sine[15382]=-19;
sine[15383]=-19;
sine[15384]=-19;
sine[15385]=-19;
sine[15386]=-19;
sine[15387]=-19;
sine[15388]=-19;
sine[15389]=-19;
sine[15390]=-19;
sine[15391]=-19;
sine[15392]=-19;
sine[15393]=-19;
sine[15394]=-19;
sine[15395]=-19;
sine[15396]=-19;
sine[15397]=-19;
sine[15398]=-19;
sine[15399]=-19;
sine[15400]=-19;
sine[15401]=-19;
sine[15402]=-20;
sine[15403]=-20;
sine[15404]=-20;
sine[15405]=-20;
sine[15406]=-20;
sine[15407]=-20;
sine[15408]=-20;
sine[15409]=-20;
sine[15410]=-20;
sine[15411]=-20;
sine[15412]=-20;
sine[15413]=-20;
sine[15414]=-20;
sine[15415]=-20;
sine[15416]=-20;
sine[15417]=-20;
sine[15418]=-20;
sine[15419]=-20;
sine[15420]=-20;
sine[15421]=-20;
sine[15422]=-20;
sine[15423]=-21;
sine[15424]=-21;
sine[15425]=-21;
sine[15426]=-21;
sine[15427]=-21;
sine[15428]=-21;
sine[15429]=-21;
sine[15430]=-21;
sine[15431]=-21;
sine[15432]=-21;
sine[15433]=-21;
sine[15434]=-21;
sine[15435]=-21;
sine[15436]=-21;
sine[15437]=-21;
sine[15438]=-21;
sine[15439]=-21;
sine[15440]=-21;
sine[15441]=-21;
sine[15442]=-21;
sine[15443]=-21;
sine[15444]=-22;
sine[15445]=-22;
sine[15446]=-22;
sine[15447]=-22;
sine[15448]=-22;
sine[15449]=-22;
sine[15450]=-22;
sine[15451]=-22;
sine[15452]=-22;
sine[15453]=-22;
sine[15454]=-22;
sine[15455]=-22;
sine[15456]=-22;
sine[15457]=-22;
sine[15458]=-22;
sine[15459]=-22;
sine[15460]=-22;
sine[15461]=-22;
sine[15462]=-22;
sine[15463]=-22;
sine[15464]=-22;
sine[15465]=-23;
sine[15466]=-23;
sine[15467]=-23;
sine[15468]=-23;
sine[15469]=-23;
sine[15470]=-23;
sine[15471]=-23;
sine[15472]=-23;
sine[15473]=-23;
sine[15474]=-23;
sine[15475]=-23;
sine[15476]=-23;
sine[15477]=-23;
sine[15478]=-23;
sine[15479]=-23;
sine[15480]=-23;
sine[15481]=-23;
sine[15482]=-23;
sine[15483]=-23;
sine[15484]=-23;
sine[15485]=-23;
sine[15486]=-23;
sine[15487]=-24;
sine[15488]=-24;
sine[15489]=-24;
sine[15490]=-24;
sine[15491]=-24;
sine[15492]=-24;
sine[15493]=-24;
sine[15494]=-24;
sine[15495]=-24;
sine[15496]=-24;
sine[15497]=-24;
sine[15498]=-24;
sine[15499]=-24;
sine[15500]=-24;
sine[15501]=-24;
sine[15502]=-24;
sine[15503]=-24;
sine[15504]=-24;
sine[15505]=-24;
sine[15506]=-24;
sine[15507]=-24;
sine[15508]=-25;
sine[15509]=-25;
sine[15510]=-25;
sine[15511]=-25;
sine[15512]=-25;
sine[15513]=-25;
sine[15514]=-25;
sine[15515]=-25;
sine[15516]=-25;
sine[15517]=-25;
sine[15518]=-25;
sine[15519]=-25;
sine[15520]=-25;
sine[15521]=-25;
sine[15522]=-25;
sine[15523]=-25;
sine[15524]=-25;
sine[15525]=-25;
sine[15526]=-25;
sine[15527]=-25;
sine[15528]=-25;
sine[15529]=-25;
sine[15530]=-26;
sine[15531]=-26;
sine[15532]=-26;
sine[15533]=-26;
sine[15534]=-26;
sine[15535]=-26;
sine[15536]=-26;
sine[15537]=-26;
sine[15538]=-26;
sine[15539]=-26;
sine[15540]=-26;
sine[15541]=-26;
sine[15542]=-26;
sine[15543]=-26;
sine[15544]=-26;
sine[15545]=-26;
sine[15546]=-26;
sine[15547]=-26;
sine[15548]=-26;
sine[15549]=-26;
sine[15550]=-26;
sine[15551]=-27;
sine[15552]=-27;
sine[15553]=-27;
sine[15554]=-27;
sine[15555]=-27;
sine[15556]=-27;
sine[15557]=-27;
sine[15558]=-27;
sine[15559]=-27;
sine[15560]=-27;
sine[15561]=-27;
sine[15562]=-27;
sine[15563]=-27;
sine[15564]=-27;
sine[15565]=-27;
sine[15566]=-27;
sine[15567]=-27;
sine[15568]=-27;
sine[15569]=-27;
sine[15570]=-27;
sine[15571]=-27;
sine[15572]=-27;
sine[15573]=-28;
sine[15574]=-28;
sine[15575]=-28;
sine[15576]=-28;
sine[15577]=-28;
sine[15578]=-28;
sine[15579]=-28;
sine[15580]=-28;
sine[15581]=-28;
sine[15582]=-28;
sine[15583]=-28;
sine[15584]=-28;
sine[15585]=-28;
sine[15586]=-28;
sine[15587]=-28;
sine[15588]=-28;
sine[15589]=-28;
sine[15590]=-28;
sine[15591]=-28;
sine[15592]=-28;
sine[15593]=-28;
sine[15594]=-28;
sine[15595]=-29;
sine[15596]=-29;
sine[15597]=-29;
sine[15598]=-29;
sine[15599]=-29;
sine[15600]=-29;
sine[15601]=-29;
sine[15602]=-29;
sine[15603]=-29;
sine[15604]=-29;
sine[15605]=-29;
sine[15606]=-29;
sine[15607]=-29;
sine[15608]=-29;
sine[15609]=-29;
sine[15610]=-29;
sine[15611]=-29;
sine[15612]=-29;
sine[15613]=-29;
sine[15614]=-29;
sine[15615]=-29;
sine[15616]=-29;
sine[15617]=-30;
sine[15618]=-30;
sine[15619]=-30;
sine[15620]=-30;
sine[15621]=-30;
sine[15622]=-30;
sine[15623]=-30;
sine[15624]=-30;
sine[15625]=-30;
sine[15626]=-30;
sine[15627]=-30;
sine[15628]=-30;
sine[15629]=-30;
sine[15630]=-30;
sine[15631]=-30;
sine[15632]=-30;
sine[15633]=-30;
sine[15634]=-30;
sine[15635]=-30;
sine[15636]=-30;
sine[15637]=-30;
sine[15638]=-30;
sine[15639]=-31;
sine[15640]=-31;
sine[15641]=-31;
sine[15642]=-31;
sine[15643]=-31;
sine[15644]=-31;
sine[15645]=-31;
sine[15646]=-31;
sine[15647]=-31;
sine[15648]=-31;
sine[15649]=-31;
sine[15650]=-31;
sine[15651]=-31;
sine[15652]=-31;
sine[15653]=-31;
sine[15654]=-31;
sine[15655]=-31;
sine[15656]=-31;
sine[15657]=-31;
sine[15658]=-31;
sine[15659]=-31;
sine[15660]=-31;
sine[15661]=-32;
sine[15662]=-32;
sine[15663]=-32;
sine[15664]=-32;
sine[15665]=-32;
sine[15666]=-32;
sine[15667]=-32;
sine[15668]=-32;
sine[15669]=-32;
sine[15670]=-32;
sine[15671]=-32;
sine[15672]=-32;
sine[15673]=-32;
sine[15674]=-32;
sine[15675]=-32;
sine[15676]=-32;
sine[15677]=-32;
sine[15678]=-32;
sine[15679]=-32;
sine[15680]=-32;
sine[15681]=-32;
sine[15682]=-32;
sine[15683]=-33;
sine[15684]=-33;
sine[15685]=-33;
sine[15686]=-33;
sine[15687]=-33;
sine[15688]=-33;
sine[15689]=-33;
sine[15690]=-33;
sine[15691]=-33;
sine[15692]=-33;
sine[15693]=-33;
sine[15694]=-33;
sine[15695]=-33;
sine[15696]=-33;
sine[15697]=-33;
sine[15698]=-33;
sine[15699]=-33;
sine[15700]=-33;
sine[15701]=-33;
sine[15702]=-33;
sine[15703]=-33;
sine[15704]=-33;
sine[15705]=-33;
sine[15706]=-34;
sine[15707]=-34;
sine[15708]=-34;
sine[15709]=-34;
sine[15710]=-34;
sine[15711]=-34;
sine[15712]=-34;
sine[15713]=-34;
sine[15714]=-34;
sine[15715]=-34;
sine[15716]=-34;
sine[15717]=-34;
sine[15718]=-34;
sine[15719]=-34;
sine[15720]=-34;
sine[15721]=-34;
sine[15722]=-34;
sine[15723]=-34;
sine[15724]=-34;
sine[15725]=-34;
sine[15726]=-34;
sine[15727]=-34;
sine[15728]=-35;
sine[15729]=-35;
sine[15730]=-35;
sine[15731]=-35;
sine[15732]=-35;
sine[15733]=-35;
sine[15734]=-35;
sine[15735]=-35;
sine[15736]=-35;
sine[15737]=-35;
sine[15738]=-35;
sine[15739]=-35;
sine[15740]=-35;
sine[15741]=-35;
sine[15742]=-35;
sine[15743]=-35;
sine[15744]=-35;
sine[15745]=-35;
sine[15746]=-35;
sine[15747]=-35;
sine[15748]=-35;
sine[15749]=-35;
sine[15750]=-35;
sine[15751]=-36;
sine[15752]=-36;
sine[15753]=-36;
sine[15754]=-36;
sine[15755]=-36;
sine[15756]=-36;
sine[15757]=-36;
sine[15758]=-36;
sine[15759]=-36;
sine[15760]=-36;
sine[15761]=-36;
sine[15762]=-36;
sine[15763]=-36;
sine[15764]=-36;
sine[15765]=-36;
sine[15766]=-36;
sine[15767]=-36;
sine[15768]=-36;
sine[15769]=-36;
sine[15770]=-36;
sine[15771]=-36;
sine[15772]=-36;
sine[15773]=-36;
sine[15774]=-37;
sine[15775]=-37;
sine[15776]=-37;
sine[15777]=-37;
sine[15778]=-37;
sine[15779]=-37;
sine[15780]=-37;
sine[15781]=-37;
sine[15782]=-37;
sine[15783]=-37;
sine[15784]=-37;
sine[15785]=-37;
sine[15786]=-37;
sine[15787]=-37;
sine[15788]=-37;
sine[15789]=-37;
sine[15790]=-37;
sine[15791]=-37;
sine[15792]=-37;
sine[15793]=-37;
sine[15794]=-37;
sine[15795]=-37;
sine[15796]=-37;
sine[15797]=-38;
sine[15798]=-38;
sine[15799]=-38;
sine[15800]=-38;
sine[15801]=-38;
sine[15802]=-38;
sine[15803]=-38;
sine[15804]=-38;
sine[15805]=-38;
sine[15806]=-38;
sine[15807]=-38;
sine[15808]=-38;
sine[15809]=-38;
sine[15810]=-38;
sine[15811]=-38;
sine[15812]=-38;
sine[15813]=-38;
sine[15814]=-38;
sine[15815]=-38;
sine[15816]=-38;
sine[15817]=-38;
sine[15818]=-38;
sine[15819]=-38;
sine[15820]=-38;
sine[15821]=-39;
sine[15822]=-39;
sine[15823]=-39;
sine[15824]=-39;
sine[15825]=-39;
sine[15826]=-39;
sine[15827]=-39;
sine[15828]=-39;
sine[15829]=-39;
sine[15830]=-39;
sine[15831]=-39;
sine[15832]=-39;
sine[15833]=-39;
sine[15834]=-39;
sine[15835]=-39;
sine[15836]=-39;
sine[15837]=-39;
sine[15838]=-39;
sine[15839]=-39;
sine[15840]=-39;
sine[15841]=-39;
sine[15842]=-39;
sine[15843]=-39;
sine[15844]=-40;
sine[15845]=-40;
sine[15846]=-40;
sine[15847]=-40;
sine[15848]=-40;
sine[15849]=-40;
sine[15850]=-40;
sine[15851]=-40;
sine[15852]=-40;
sine[15853]=-40;
sine[15854]=-40;
sine[15855]=-40;
sine[15856]=-40;
sine[15857]=-40;
sine[15858]=-40;
sine[15859]=-40;
sine[15860]=-40;
sine[15861]=-40;
sine[15862]=-40;
sine[15863]=-40;
sine[15864]=-40;
sine[15865]=-40;
sine[15866]=-40;
sine[15867]=-40;
sine[15868]=-41;
sine[15869]=-41;
sine[15870]=-41;
sine[15871]=-41;
sine[15872]=-41;
sine[15873]=-41;
sine[15874]=-41;
sine[15875]=-41;
sine[15876]=-41;
sine[15877]=-41;
sine[15878]=-41;
sine[15879]=-41;
sine[15880]=-41;
sine[15881]=-41;
sine[15882]=-41;
sine[15883]=-41;
sine[15884]=-41;
sine[15885]=-41;
sine[15886]=-41;
sine[15887]=-41;
sine[15888]=-41;
sine[15889]=-41;
sine[15890]=-41;
sine[15891]=-41;
sine[15892]=-42;
sine[15893]=-42;
sine[15894]=-42;
sine[15895]=-42;
sine[15896]=-42;
sine[15897]=-42;
sine[15898]=-42;
sine[15899]=-42;
sine[15900]=-42;
sine[15901]=-42;
sine[15902]=-42;
sine[15903]=-42;
sine[15904]=-42;
sine[15905]=-42;
sine[15906]=-42;
sine[15907]=-42;
sine[15908]=-42;
sine[15909]=-42;
sine[15910]=-42;
sine[15911]=-42;
sine[15912]=-42;
sine[15913]=-42;
sine[15914]=-42;
sine[15915]=-42;
sine[15916]=-43;
sine[15917]=-43;
sine[15918]=-43;
sine[15919]=-43;
sine[15920]=-43;
sine[15921]=-43;
sine[15922]=-43;
sine[15923]=-43;
sine[15924]=-43;
sine[15925]=-43;
sine[15926]=-43;
sine[15927]=-43;
sine[15928]=-43;
sine[15929]=-43;
sine[15930]=-43;
sine[15931]=-43;
sine[15932]=-43;
sine[15933]=-43;
sine[15934]=-43;
sine[15935]=-43;
sine[15936]=-43;
sine[15937]=-43;
sine[15938]=-43;
sine[15939]=-43;
sine[15940]=-44;
sine[15941]=-44;
sine[15942]=-44;
sine[15943]=-44;
sine[15944]=-44;
sine[15945]=-44;
sine[15946]=-44;
sine[15947]=-44;
sine[15948]=-44;
sine[15949]=-44;
sine[15950]=-44;
sine[15951]=-44;
sine[15952]=-44;
sine[15953]=-44;
sine[15954]=-44;
sine[15955]=-44;
sine[15956]=-44;
sine[15957]=-44;
sine[15958]=-44;
sine[15959]=-44;
sine[15960]=-44;
sine[15961]=-44;
sine[15962]=-44;
sine[15963]=-44;
sine[15964]=-44;
sine[15965]=-45;
sine[15966]=-45;
sine[15967]=-45;
sine[15968]=-45;
sine[15969]=-45;
sine[15970]=-45;
sine[15971]=-45;
sine[15972]=-45;
sine[15973]=-45;
sine[15974]=-45;
sine[15975]=-45;
sine[15976]=-45;
sine[15977]=-45;
sine[15978]=-45;
sine[15979]=-45;
sine[15980]=-45;
sine[15981]=-45;
sine[15982]=-45;
sine[15983]=-45;
sine[15984]=-45;
sine[15985]=-45;
sine[15986]=-45;
sine[15987]=-45;
sine[15988]=-45;
sine[15989]=-45;
sine[15990]=-46;
sine[15991]=-46;
sine[15992]=-46;
sine[15993]=-46;
sine[15994]=-46;
sine[15995]=-46;
sine[15996]=-46;
sine[15997]=-46;
sine[15998]=-46;
sine[15999]=-46;
sine[16000]=-46;
sine[16001]=-46;
sine[16002]=-46;
sine[16003]=-46;
sine[16004]=-46;
sine[16005]=-46;
sine[16006]=-46;
sine[16007]=-46;
sine[16008]=-46;
sine[16009]=-46;
sine[16010]=-46;
sine[16011]=-46;
sine[16012]=-46;
sine[16013]=-46;
sine[16014]=-46;
sine[16015]=-47;
sine[16016]=-47;
sine[16017]=-47;
sine[16018]=-47;
sine[16019]=-47;
sine[16020]=-47;
sine[16021]=-47;
sine[16022]=-47;
sine[16023]=-47;
sine[16024]=-47;
sine[16025]=-47;
sine[16026]=-47;
sine[16027]=-47;
sine[16028]=-47;
sine[16029]=-47;
sine[16030]=-47;
sine[16031]=-47;
sine[16032]=-47;
sine[16033]=-47;
sine[16034]=-47;
sine[16035]=-47;
sine[16036]=-47;
sine[16037]=-47;
sine[16038]=-47;
sine[16039]=-47;
sine[16040]=-47;
sine[16041]=-48;
sine[16042]=-48;
sine[16043]=-48;
sine[16044]=-48;
sine[16045]=-48;
sine[16046]=-48;
sine[16047]=-48;
sine[16048]=-48;
sine[16049]=-48;
sine[16050]=-48;
sine[16051]=-48;
sine[16052]=-48;
sine[16053]=-48;
sine[16054]=-48;
sine[16055]=-48;
sine[16056]=-48;
sine[16057]=-48;
sine[16058]=-48;
sine[16059]=-48;
sine[16060]=-48;
sine[16061]=-48;
sine[16062]=-48;
sine[16063]=-48;
sine[16064]=-48;
sine[16065]=-48;
sine[16066]=-49;
sine[16067]=-49;
sine[16068]=-49;
sine[16069]=-49;
sine[16070]=-49;
sine[16071]=-49;
sine[16072]=-49;
sine[16073]=-49;
sine[16074]=-49;
sine[16075]=-49;
sine[16076]=-49;
sine[16077]=-49;
sine[16078]=-49;
sine[16079]=-49;
sine[16080]=-49;
sine[16081]=-49;
sine[16082]=-49;
sine[16083]=-49;
sine[16084]=-49;
sine[16085]=-49;
sine[16086]=-49;
sine[16087]=-49;
sine[16088]=-49;
sine[16089]=-49;
sine[16090]=-49;
sine[16091]=-49;
sine[16092]=-49;
sine[16093]=-50;
sine[16094]=-50;
sine[16095]=-50;
sine[16096]=-50;
sine[16097]=-50;
sine[16098]=-50;
sine[16099]=-50;
sine[16100]=-50;
sine[16101]=-50;
sine[16102]=-50;
sine[16103]=-50;
sine[16104]=-50;
sine[16105]=-50;
sine[16106]=-50;
sine[16107]=-50;
sine[16108]=-50;
sine[16109]=-50;
sine[16110]=-50;
sine[16111]=-50;
sine[16112]=-50;
sine[16113]=-50;
sine[16114]=-50;
sine[16115]=-50;
sine[16116]=-50;
sine[16117]=-50;
sine[16118]=-50;
sine[16119]=-51;
sine[16120]=-51;
sine[16121]=-51;
sine[16122]=-51;
sine[16123]=-51;
sine[16124]=-51;
sine[16125]=-51;
sine[16126]=-51;
sine[16127]=-51;
sine[16128]=-51;
sine[16129]=-51;
sine[16130]=-51;
sine[16131]=-51;
sine[16132]=-51;
sine[16133]=-51;
sine[16134]=-51;
sine[16135]=-51;
sine[16136]=-51;
sine[16137]=-51;
sine[16138]=-51;
sine[16139]=-51;
sine[16140]=-51;
sine[16141]=-51;
sine[16142]=-51;
sine[16143]=-51;
sine[16144]=-51;
sine[16145]=-51;
sine[16146]=-52;
sine[16147]=-52;
sine[16148]=-52;
sine[16149]=-52;
sine[16150]=-52;
sine[16151]=-52;
sine[16152]=-52;
sine[16153]=-52;
sine[16154]=-52;
sine[16155]=-52;
sine[16156]=-52;
sine[16157]=-52;
sine[16158]=-52;
sine[16159]=-52;
sine[16160]=-52;
sine[16161]=-52;
sine[16162]=-52;
sine[16163]=-52;
sine[16164]=-52;
sine[16165]=-52;
sine[16166]=-52;
sine[16167]=-52;
sine[16168]=-52;
sine[16169]=-52;
sine[16170]=-52;
sine[16171]=-52;
sine[16172]=-52;
sine[16173]=-53;
sine[16174]=-53;
sine[16175]=-53;
sine[16176]=-53;
sine[16177]=-53;
sine[16178]=-53;
sine[16179]=-53;
sine[16180]=-53;
sine[16181]=-53;
sine[16182]=-53;
sine[16183]=-53;
sine[16184]=-53;
sine[16185]=-53;
sine[16186]=-53;
sine[16187]=-53;
sine[16188]=-53;
sine[16189]=-53;
sine[16190]=-53;
sine[16191]=-53;
sine[16192]=-53;
sine[16193]=-53;
sine[16194]=-53;
sine[16195]=-53;
sine[16196]=-53;
sine[16197]=-53;
sine[16198]=-53;
sine[16199]=-53;
sine[16200]=-53;
sine[16201]=-54;
sine[16202]=-54;
sine[16203]=-54;
sine[16204]=-54;
sine[16205]=-54;
sine[16206]=-54;
sine[16207]=-54;
sine[16208]=-54;
sine[16209]=-54;
sine[16210]=-54;
sine[16211]=-54;
sine[16212]=-54;
sine[16213]=-54;
sine[16214]=-54;
sine[16215]=-54;
sine[16216]=-54;
sine[16217]=-54;
sine[16218]=-54;
sine[16219]=-54;
sine[16220]=-54;
sine[16221]=-54;
sine[16222]=-54;
sine[16223]=-54;
sine[16224]=-54;
sine[16225]=-54;
sine[16226]=-54;
sine[16227]=-54;
sine[16228]=-54;
sine[16229]=-55;
sine[16230]=-55;
sine[16231]=-55;
sine[16232]=-55;
sine[16233]=-55;
sine[16234]=-55;
sine[16235]=-55;
sine[16236]=-55;
sine[16237]=-55;
sine[16238]=-55;
sine[16239]=-55;
sine[16240]=-55;
sine[16241]=-55;
sine[16242]=-55;
sine[16243]=-55;
sine[16244]=-55;
sine[16245]=-55;
sine[16246]=-55;
sine[16247]=-55;
sine[16248]=-55;
sine[16249]=-55;
sine[16250]=-55;
sine[16251]=-55;
sine[16252]=-55;
sine[16253]=-55;
sine[16254]=-55;
sine[16255]=-55;
sine[16256]=-55;
sine[16257]=-55;
sine[16258]=-56;
sine[16259]=-56;
sine[16260]=-56;
sine[16261]=-56;
sine[16262]=-56;
sine[16263]=-56;
sine[16264]=-56;
sine[16265]=-56;
sine[16266]=-56;
sine[16267]=-56;
sine[16268]=-56;
sine[16269]=-56;
sine[16270]=-56;
sine[16271]=-56;
sine[16272]=-56;
sine[16273]=-56;
sine[16274]=-56;
sine[16275]=-56;
sine[16276]=-56;
sine[16277]=-56;
sine[16278]=-56;
sine[16279]=-56;
sine[16280]=-56;
sine[16281]=-56;
sine[16282]=-56;
sine[16283]=-56;
sine[16284]=-56;
sine[16285]=-56;
sine[16286]=-56;
sine[16287]=-57;
sine[16288]=-57;
sine[16289]=-57;
sine[16290]=-57;
sine[16291]=-57;
sine[16292]=-57;
sine[16293]=-57;
sine[16294]=-57;
sine[16295]=-57;
sine[16296]=-57;
sine[16297]=-57;
sine[16298]=-57;
sine[16299]=-57;
sine[16300]=-57;
sine[16301]=-57;
sine[16302]=-57;
sine[16303]=-57;
sine[16304]=-57;
sine[16305]=-57;
sine[16306]=-57;
sine[16307]=-57;
sine[16308]=-57;
sine[16309]=-57;
sine[16310]=-57;
sine[16311]=-57;
sine[16312]=-57;
sine[16313]=-57;
sine[16314]=-57;
sine[16315]=-57;
sine[16316]=-57;
sine[16317]=-58;
sine[16318]=-58;
sine[16319]=-58;
sine[16320]=-58;
sine[16321]=-58;
sine[16322]=-58;
sine[16323]=-58;
sine[16324]=-58;
sine[16325]=-58;
sine[16326]=-58;
sine[16327]=-58;
sine[16328]=-58;
sine[16329]=-58;
sine[16330]=-58;
sine[16331]=-58;
sine[16332]=-58;
sine[16333]=-58;
sine[16334]=-58;
sine[16335]=-58;
sine[16336]=-58;
sine[16337]=-58;
sine[16338]=-58;
sine[16339]=-58;
sine[16340]=-58;
sine[16341]=-58;
sine[16342]=-58;
sine[16343]=-58;
sine[16344]=-58;
sine[16345]=-58;
sine[16346]=-58;
sine[16347]=-59;
sine[16348]=-59;
sine[16349]=-59;
sine[16350]=-59;
sine[16351]=-59;
sine[16352]=-59;
sine[16353]=-59;
sine[16354]=-59;
sine[16355]=-59;
sine[16356]=-59;
sine[16357]=-59;
sine[16358]=-59;
sine[16359]=-59;
sine[16360]=-59;
sine[16361]=-59;
sine[16362]=-59;
sine[16363]=-59;
sine[16364]=-59;
sine[16365]=-59;
sine[16366]=-59;
sine[16367]=-59;
sine[16368]=-59;
sine[16369]=-59;
sine[16370]=-59;
sine[16371]=-59;
sine[16372]=-59;
sine[16373]=-59;
sine[16374]=-59;
sine[16375]=-59;
sine[16376]=-59;
sine[16377]=-59;
sine[16378]=-60;
sine[16379]=-60;
sine[16380]=-60;
sine[16381]=-60;
sine[16382]=-60;
sine[16383]=-60;
sine[16384]=-60;
sine[16385]=-60;
sine[16386]=-60;
sine[16387]=-60;
sine[16388]=-60;
sine[16389]=-60;
sine[16390]=-60;
sine[16391]=-60;
sine[16392]=-60;
sine[16393]=-60;
sine[16394]=-60;
sine[16395]=-60;
sine[16396]=-60;
sine[16397]=-60;
sine[16398]=-60;
sine[16399]=-60;
sine[16400]=-60;
sine[16401]=-60;
sine[16402]=-60;
sine[16403]=-60;
sine[16404]=-60;
sine[16405]=-60;
sine[16406]=-60;
sine[16407]=-60;
sine[16408]=-60;
sine[16409]=-60;
sine[16410]=-61;
sine[16411]=-61;
sine[16412]=-61;
sine[16413]=-61;
sine[16414]=-61;
sine[16415]=-61;
sine[16416]=-61;
sine[16417]=-61;
sine[16418]=-61;
sine[16419]=-61;
sine[16420]=-61;
sine[16421]=-61;
sine[16422]=-61;
sine[16423]=-61;
sine[16424]=-61;
sine[16425]=-61;
sine[16426]=-61;
sine[16427]=-61;
sine[16428]=-61;
sine[16429]=-61;
sine[16430]=-61;
sine[16431]=-61;
sine[16432]=-61;
sine[16433]=-61;
sine[16434]=-61;
sine[16435]=-61;
sine[16436]=-61;
sine[16437]=-61;
sine[16438]=-61;
sine[16439]=-61;
sine[16440]=-61;
sine[16441]=-61;
sine[16442]=-61;
sine[16443]=-62;
sine[16444]=-62;
sine[16445]=-62;
sine[16446]=-62;
sine[16447]=-62;
sine[16448]=-62;
sine[16449]=-62;
sine[16450]=-62;
sine[16451]=-62;
sine[16452]=-62;
sine[16453]=-62;
sine[16454]=-62;
sine[16455]=-62;
sine[16456]=-62;
sine[16457]=-62;
sine[16458]=-62;
sine[16459]=-62;
sine[16460]=-62;
sine[16461]=-62;
sine[16462]=-62;
sine[16463]=-62;
sine[16464]=-62;
sine[16465]=-62;
sine[16466]=-62;
sine[16467]=-62;
sine[16468]=-62;
sine[16469]=-62;
sine[16470]=-62;
sine[16471]=-62;
sine[16472]=-62;
sine[16473]=-62;
sine[16474]=-62;
sine[16475]=-62;
sine[16476]=-63;
sine[16477]=-63;
sine[16478]=-63;
sine[16479]=-63;
sine[16480]=-63;
sine[16481]=-63;
sine[16482]=-63;
sine[16483]=-63;
sine[16484]=-63;
sine[16485]=-63;
sine[16486]=-63;
sine[16487]=-63;
sine[16488]=-63;
sine[16489]=-63;
sine[16490]=-63;
sine[16491]=-63;
sine[16492]=-63;
sine[16493]=-63;
sine[16494]=-63;
sine[16495]=-63;
sine[16496]=-63;
sine[16497]=-63;
sine[16498]=-63;
sine[16499]=-63;
sine[16500]=-63;
sine[16501]=-63;
sine[16502]=-63;
sine[16503]=-63;
sine[16504]=-63;
sine[16505]=-63;
sine[16506]=-63;
sine[16507]=-63;
sine[16508]=-63;
sine[16509]=-63;
sine[16510]=-63;
sine[16511]=-64;
sine[16512]=-64;
sine[16513]=-64;
sine[16514]=-64;
sine[16515]=-64;
sine[16516]=-64;
sine[16517]=-64;
sine[16518]=-64;
sine[16519]=-64;
sine[16520]=-64;
sine[16521]=-64;
sine[16522]=-64;
sine[16523]=-64;
sine[16524]=-64;
sine[16525]=-64;
sine[16526]=-64;
sine[16527]=-64;
sine[16528]=-64;
sine[16529]=-64;
sine[16530]=-64;
sine[16531]=-64;
sine[16532]=-64;
sine[16533]=-64;
sine[16534]=-64;
sine[16535]=-64;
sine[16536]=-64;
sine[16537]=-64;
sine[16538]=-64;
sine[16539]=-64;
sine[16540]=-64;
sine[16541]=-64;
sine[16542]=-64;
sine[16543]=-64;
sine[16544]=-64;
sine[16545]=-64;
sine[16546]=-65;
sine[16547]=-65;
sine[16548]=-65;
sine[16549]=-65;
sine[16550]=-65;
sine[16551]=-65;
sine[16552]=-65;
sine[16553]=-65;
sine[16554]=-65;
sine[16555]=-65;
sine[16556]=-65;
sine[16557]=-65;
sine[16558]=-65;
sine[16559]=-65;
sine[16560]=-65;
sine[16561]=-65;
sine[16562]=-65;
sine[16563]=-65;
sine[16564]=-65;
sine[16565]=-65;
sine[16566]=-65;
sine[16567]=-65;
sine[16568]=-65;
sine[16569]=-65;
sine[16570]=-65;
sine[16571]=-65;
sine[16572]=-65;
sine[16573]=-65;
sine[16574]=-65;
sine[16575]=-65;
sine[16576]=-65;
sine[16577]=-65;
sine[16578]=-65;
sine[16579]=-65;
sine[16580]=-65;
sine[16581]=-65;
sine[16582]=-65;
sine[16583]=-66;
sine[16584]=-66;
sine[16585]=-66;
sine[16586]=-66;
sine[16587]=-66;
sine[16588]=-66;
sine[16589]=-66;
sine[16590]=-66;
sine[16591]=-66;
sine[16592]=-66;
sine[16593]=-66;
sine[16594]=-66;
sine[16595]=-66;
sine[16596]=-66;
sine[16597]=-66;
sine[16598]=-66;
sine[16599]=-66;
sine[16600]=-66;
sine[16601]=-66;
sine[16602]=-66;
sine[16603]=-66;
sine[16604]=-66;
sine[16605]=-66;
sine[16606]=-66;
sine[16607]=-66;
sine[16608]=-66;
sine[16609]=-66;
sine[16610]=-66;
sine[16611]=-66;
sine[16612]=-66;
sine[16613]=-66;
sine[16614]=-66;
sine[16615]=-66;
sine[16616]=-66;
sine[16617]=-66;
sine[16618]=-66;
sine[16619]=-66;
sine[16620]=-66;
sine[16621]=-67;
sine[16622]=-67;
sine[16623]=-67;
sine[16624]=-67;
sine[16625]=-67;
sine[16626]=-67;
sine[16627]=-67;
sine[16628]=-67;
sine[16629]=-67;
sine[16630]=-67;
sine[16631]=-67;
sine[16632]=-67;
sine[16633]=-67;
sine[16634]=-67;
sine[16635]=-67;
sine[16636]=-67;
sine[16637]=-67;
sine[16638]=-67;
sine[16639]=-67;
sine[16640]=-67;
sine[16641]=-67;
sine[16642]=-67;
sine[16643]=-67;
sine[16644]=-67;
sine[16645]=-67;
sine[16646]=-67;
sine[16647]=-67;
sine[16648]=-67;
sine[16649]=-67;
sine[16650]=-67;
sine[16651]=-67;
sine[16652]=-67;
sine[16653]=-67;
sine[16654]=-67;
sine[16655]=-67;
sine[16656]=-67;
sine[16657]=-67;
sine[16658]=-67;
sine[16659]=-67;
sine[16660]=-67;
sine[16661]=-68;
sine[16662]=-68;
sine[16663]=-68;
sine[16664]=-68;
sine[16665]=-68;
sine[16666]=-68;
sine[16667]=-68;
sine[16668]=-68;
sine[16669]=-68;
sine[16670]=-68;
sine[16671]=-68;
sine[16672]=-68;
sine[16673]=-68;
sine[16674]=-68;
sine[16675]=-68;
sine[16676]=-68;
sine[16677]=-68;
sine[16678]=-68;
sine[16679]=-68;
sine[16680]=-68;
sine[16681]=-68;
sine[16682]=-68;
sine[16683]=-68;
sine[16684]=-68;
sine[16685]=-68;
sine[16686]=-68;
sine[16687]=-68;
sine[16688]=-68;
sine[16689]=-68;
sine[16690]=-68;
sine[16691]=-68;
sine[16692]=-68;
sine[16693]=-68;
sine[16694]=-68;
sine[16695]=-68;
sine[16696]=-68;
sine[16697]=-68;
sine[16698]=-68;
sine[16699]=-68;
sine[16700]=-68;
sine[16701]=-68;
sine[16702]=-69;
sine[16703]=-69;
sine[16704]=-69;
sine[16705]=-69;
sine[16706]=-69;
sine[16707]=-69;
sine[16708]=-69;
sine[16709]=-69;
sine[16710]=-69;
sine[16711]=-69;
sine[16712]=-69;
sine[16713]=-69;
sine[16714]=-69;
sine[16715]=-69;
sine[16716]=-69;
sine[16717]=-69;
sine[16718]=-69;
sine[16719]=-69;
sine[16720]=-69;
sine[16721]=-69;
sine[16722]=-69;
sine[16723]=-69;
sine[16724]=-69;
sine[16725]=-69;
sine[16726]=-69;
sine[16727]=-69;
sine[16728]=-69;
sine[16729]=-69;
sine[16730]=-69;
sine[16731]=-69;
sine[16732]=-69;
sine[16733]=-69;
sine[16734]=-69;
sine[16735]=-69;
sine[16736]=-69;
sine[16737]=-69;
sine[16738]=-69;
sine[16739]=-69;
sine[16740]=-69;
sine[16741]=-69;
sine[16742]=-69;
sine[16743]=-69;
sine[16744]=-69;
sine[16745]=-69;
sine[16746]=-70;
sine[16747]=-70;
sine[16748]=-70;
sine[16749]=-70;
sine[16750]=-70;
sine[16751]=-70;
sine[16752]=-70;
sine[16753]=-70;
sine[16754]=-70;
sine[16755]=-70;
sine[16756]=-70;
sine[16757]=-70;
sine[16758]=-70;
sine[16759]=-70;
sine[16760]=-70;
sine[16761]=-70;
sine[16762]=-70;
sine[16763]=-70;
sine[16764]=-70;
sine[16765]=-70;
sine[16766]=-70;
sine[16767]=-70;
sine[16768]=-70;
sine[16769]=-70;
sine[16770]=-70;
sine[16771]=-70;
sine[16772]=-70;
sine[16773]=-70;
sine[16774]=-70;
sine[16775]=-70;
sine[16776]=-70;
sine[16777]=-70;
sine[16778]=-70;
sine[16779]=-70;
sine[16780]=-70;
sine[16781]=-70;
sine[16782]=-70;
sine[16783]=-70;
sine[16784]=-70;
sine[16785]=-70;
sine[16786]=-70;
sine[16787]=-70;
sine[16788]=-70;
sine[16789]=-70;
sine[16790]=-70;
sine[16791]=-71;
sine[16792]=-71;
sine[16793]=-71;
sine[16794]=-71;
sine[16795]=-71;
sine[16796]=-71;
sine[16797]=-71;
sine[16798]=-71;
sine[16799]=-71;
sine[16800]=-71;
sine[16801]=-71;
sine[16802]=-71;
sine[16803]=-71;
sine[16804]=-71;
sine[16805]=-71;
sine[16806]=-71;
sine[16807]=-71;
sine[16808]=-71;
sine[16809]=-71;
sine[16810]=-71;
sine[16811]=-71;
sine[16812]=-71;
sine[16813]=-71;
sine[16814]=-71;
sine[16815]=-71;
sine[16816]=-71;
sine[16817]=-71;
sine[16818]=-71;
sine[16819]=-71;
sine[16820]=-71;
sine[16821]=-71;
sine[16822]=-71;
sine[16823]=-71;
sine[16824]=-71;
sine[16825]=-71;
sine[16826]=-71;
sine[16827]=-71;
sine[16828]=-71;
sine[16829]=-71;
sine[16830]=-71;
sine[16831]=-71;
sine[16832]=-71;
sine[16833]=-71;
sine[16834]=-71;
sine[16835]=-71;
sine[16836]=-71;
sine[16837]=-71;
sine[16838]=-71;
sine[16839]=-71;
sine[16840]=-72;
sine[16841]=-72;
sine[16842]=-72;
sine[16843]=-72;
sine[16844]=-72;
sine[16845]=-72;
sine[16846]=-72;
sine[16847]=-72;
sine[16848]=-72;
sine[16849]=-72;
sine[16850]=-72;
sine[16851]=-72;
sine[16852]=-72;
sine[16853]=-72;
sine[16854]=-72;
sine[16855]=-72;
sine[16856]=-72;
sine[16857]=-72;
sine[16858]=-72;
sine[16859]=-72;
sine[16860]=-72;
sine[16861]=-72;
sine[16862]=-72;
sine[16863]=-72;
sine[16864]=-72;
sine[16865]=-72;
sine[16866]=-72;
sine[16867]=-72;
sine[16868]=-72;
sine[16869]=-72;
sine[16870]=-72;
sine[16871]=-72;
sine[16872]=-72;
sine[16873]=-72;
sine[16874]=-72;
sine[16875]=-72;
sine[16876]=-72;
sine[16877]=-72;
sine[16878]=-72;
sine[16879]=-72;
sine[16880]=-72;
sine[16881]=-72;
sine[16882]=-72;
sine[16883]=-72;
sine[16884]=-72;
sine[16885]=-72;
sine[16886]=-72;
sine[16887]=-72;
sine[16888]=-72;
sine[16889]=-72;
sine[16890]=-72;
sine[16891]=-72;
sine[16892]=-72;
sine[16893]=-73;
sine[16894]=-73;
sine[16895]=-73;
sine[16896]=-73;
sine[16897]=-73;
sine[16898]=-73;
sine[16899]=-73;
sine[16900]=-73;
sine[16901]=-73;
sine[16902]=-73;
sine[16903]=-73;
sine[16904]=-73;
sine[16905]=-73;
sine[16906]=-73;
sine[16907]=-73;
sine[16908]=-73;
sine[16909]=-73;
sine[16910]=-73;
sine[16911]=-73;
sine[16912]=-73;
sine[16913]=-73;
sine[16914]=-73;
sine[16915]=-73;
sine[16916]=-73;
sine[16917]=-73;
sine[16918]=-73;
sine[16919]=-73;
sine[16920]=-73;
sine[16921]=-73;
sine[16922]=-73;
sine[16923]=-73;
sine[16924]=-73;
sine[16925]=-73;
sine[16926]=-73;
sine[16927]=-73;
sine[16928]=-73;
sine[16929]=-73;
sine[16930]=-73;
sine[16931]=-73;
sine[16932]=-73;
sine[16933]=-73;
sine[16934]=-73;
sine[16935]=-73;
sine[16936]=-73;
sine[16937]=-73;
sine[16938]=-73;
sine[16939]=-73;
sine[16940]=-73;
sine[16941]=-73;
sine[16942]=-73;
sine[16943]=-73;
sine[16944]=-73;
sine[16945]=-73;
sine[16946]=-73;
sine[16947]=-73;
sine[16948]=-73;
sine[16949]=-73;
sine[16950]=-74;
sine[16951]=-74;
sine[16952]=-74;
sine[16953]=-74;
sine[16954]=-74;
sine[16955]=-74;
sine[16956]=-74;
sine[16957]=-74;
sine[16958]=-74;
sine[16959]=-74;
sine[16960]=-74;
sine[16961]=-74;
sine[16962]=-74;
sine[16963]=-74;
sine[16964]=-74;
sine[16965]=-74;
sine[16966]=-74;
sine[16967]=-74;
sine[16968]=-74;
sine[16969]=-74;
sine[16970]=-74;
sine[16971]=-74;
sine[16972]=-74;
sine[16973]=-74;
sine[16974]=-74;
sine[16975]=-74;
sine[16976]=-74;
sine[16977]=-74;
sine[16978]=-74;
sine[16979]=-74;
sine[16980]=-74;
sine[16981]=-74;
sine[16982]=-74;
sine[16983]=-74;
sine[16984]=-74;
sine[16985]=-74;
sine[16986]=-74;
sine[16987]=-74;
sine[16988]=-74;
sine[16989]=-74;
sine[16990]=-74;
sine[16991]=-74;
sine[16992]=-74;
sine[16993]=-74;
sine[16994]=-74;
sine[16995]=-74;
sine[16996]=-74;
sine[16997]=-74;
sine[16998]=-74;
sine[16999]=-74;
sine[17000]=-74;
sine[17001]=-74;
sine[17002]=-74;
sine[17003]=-74;
sine[17004]=-74;
sine[17005]=-74;
sine[17006]=-74;
sine[17007]=-74;
sine[17008]=-74;
sine[17009]=-74;
sine[17010]=-74;
sine[17011]=-74;
sine[17012]=-74;
sine[17013]=-74;
sine[17014]=-75;
sine[17015]=-75;
sine[17016]=-75;
sine[17017]=-75;
sine[17018]=-75;
sine[17019]=-75;
sine[17020]=-75;
sine[17021]=-75;
sine[17022]=-75;
sine[17023]=-75;
sine[17024]=-75;
sine[17025]=-75;
sine[17026]=-75;
sine[17027]=-75;
sine[17028]=-75;
sine[17029]=-75;
sine[17030]=-75;
sine[17031]=-75;
sine[17032]=-75;
sine[17033]=-75;
sine[17034]=-75;
sine[17035]=-75;
sine[17036]=-75;
sine[17037]=-75;
sine[17038]=-75;
sine[17039]=-75;
sine[17040]=-75;
sine[17041]=-75;
sine[17042]=-75;
sine[17043]=-75;
sine[17044]=-75;
sine[17045]=-75;
sine[17046]=-75;
sine[17047]=-75;
sine[17048]=-75;
sine[17049]=-75;
sine[17050]=-75;
sine[17051]=-75;
sine[17052]=-75;
sine[17053]=-75;
sine[17054]=-75;
sine[17055]=-75;
sine[17056]=-75;
sine[17057]=-75;
sine[17058]=-75;
sine[17059]=-75;
sine[17060]=-75;
sine[17061]=-75;
sine[17062]=-75;
sine[17063]=-75;
sine[17064]=-75;
sine[17065]=-75;
sine[17066]=-75;
sine[17067]=-75;
sine[17068]=-75;
sine[17069]=-75;
sine[17070]=-75;
sine[17071]=-75;
sine[17072]=-75;
sine[17073]=-75;
sine[17074]=-75;
sine[17075]=-75;
sine[17076]=-75;
sine[17077]=-75;
sine[17078]=-75;
sine[17079]=-75;
sine[17080]=-75;
sine[17081]=-75;
sine[17082]=-75;
sine[17083]=-75;
sine[17084]=-75;
sine[17085]=-75;
sine[17086]=-75;
sine[17087]=-76;
sine[17088]=-76;
sine[17089]=-76;
sine[17090]=-76;
sine[17091]=-76;
sine[17092]=-76;
sine[17093]=-76;
sine[17094]=-76;
sine[17095]=-76;
sine[17096]=-76;
sine[17097]=-76;
sine[17098]=-76;
sine[17099]=-76;
sine[17100]=-76;
sine[17101]=-76;
sine[17102]=-76;
sine[17103]=-76;
sine[17104]=-76;
sine[17105]=-76;
sine[17106]=-76;
sine[17107]=-76;
sine[17108]=-76;
sine[17109]=-76;
sine[17110]=-76;
sine[17111]=-76;
sine[17112]=-76;
sine[17113]=-76;
sine[17114]=-76;
sine[17115]=-76;
sine[17116]=-76;
sine[17117]=-76;
sine[17118]=-76;
sine[17119]=-76;
sine[17120]=-76;
sine[17121]=-76;
sine[17122]=-76;
sine[17123]=-76;
sine[17124]=-76;
sine[17125]=-76;
sine[17126]=-76;
sine[17127]=-76;
sine[17128]=-76;
sine[17129]=-76;
sine[17130]=-76;
sine[17131]=-76;
sine[17132]=-76;
sine[17133]=-76;
sine[17134]=-76;
sine[17135]=-76;
sine[17136]=-76;
sine[17137]=-76;
sine[17138]=-76;
sine[17139]=-76;
sine[17140]=-76;
sine[17141]=-76;
sine[17142]=-76;
sine[17143]=-76;
sine[17144]=-76;
sine[17145]=-76;
sine[17146]=-76;
sine[17147]=-76;
sine[17148]=-76;
sine[17149]=-76;
sine[17150]=-76;
sine[17151]=-76;
sine[17152]=-76;
sine[17153]=-76;
sine[17154]=-76;
sine[17155]=-76;
sine[17156]=-76;
sine[17157]=-76;
sine[17158]=-76;
sine[17159]=-76;
sine[17160]=-76;
sine[17161]=-76;
sine[17162]=-76;
sine[17163]=-76;
sine[17164]=-76;
sine[17165]=-76;
sine[17166]=-76;
sine[17167]=-76;
sine[17168]=-76;
sine[17169]=-76;
sine[17170]=-76;
sine[17171]=-76;
sine[17172]=-76;
sine[17173]=-76;
sine[17174]=-76;
sine[17175]=-77;
sine[17176]=-77;
sine[17177]=-77;
sine[17178]=-77;
sine[17179]=-77;
sine[17180]=-77;
sine[17181]=-77;
sine[17182]=-77;
sine[17183]=-77;
sine[17184]=-77;
sine[17185]=-77;
sine[17186]=-77;
sine[17187]=-77;
sine[17188]=-77;
sine[17189]=-77;
sine[17190]=-77;
sine[17191]=-77;
sine[17192]=-77;
sine[17193]=-77;
sine[17194]=-77;
sine[17195]=-77;
sine[17196]=-77;
sine[17197]=-77;
sine[17198]=-77;
sine[17199]=-77;
sine[17200]=-77;
sine[17201]=-77;
sine[17202]=-77;
sine[17203]=-77;
sine[17204]=-77;
sine[17205]=-77;
sine[17206]=-77;
sine[17207]=-77;
sine[17208]=-77;
sine[17209]=-77;
sine[17210]=-77;
sine[17211]=-77;
sine[17212]=-77;
sine[17213]=-77;
sine[17214]=-77;
sine[17215]=-77;
sine[17216]=-77;
sine[17217]=-77;
sine[17218]=-77;
sine[17219]=-77;
sine[17220]=-77;
sine[17221]=-77;
sine[17222]=-77;
sine[17223]=-77;
sine[17224]=-77;
sine[17225]=-77;
sine[17226]=-77;
sine[17227]=-77;
sine[17228]=-77;
sine[17229]=-77;
sine[17230]=-77;
sine[17231]=-77;
sine[17232]=-77;
sine[17233]=-77;
sine[17234]=-77;
sine[17235]=-77;
sine[17236]=-77;
sine[17237]=-77;
sine[17238]=-77;
sine[17239]=-77;
sine[17240]=-77;
sine[17241]=-77;
sine[17242]=-77;
sine[17243]=-77;
sine[17244]=-77;
sine[17245]=-77;
sine[17246]=-77;
sine[17247]=-77;
sine[17248]=-77;
sine[17249]=-77;
sine[17250]=-77;
sine[17251]=-77;
sine[17252]=-77;
sine[17253]=-77;
sine[17254]=-77;
sine[17255]=-77;
sine[17256]=-77;
sine[17257]=-77;
sine[17258]=-77;
sine[17259]=-77;
sine[17260]=-77;
sine[17261]=-77;
sine[17262]=-77;
sine[17263]=-77;
sine[17264]=-77;
sine[17265]=-77;
sine[17266]=-77;
sine[17267]=-77;
sine[17268]=-77;
sine[17269]=-77;
sine[17270]=-77;
sine[17271]=-77;
sine[17272]=-77;
sine[17273]=-77;
sine[17274]=-77;
sine[17275]=-77;
sine[17276]=-77;
sine[17277]=-77;
sine[17278]=-77;
sine[17279]=-77;
sine[17280]=-77;
sine[17281]=-77;
sine[17282]=-77;
sine[17283]=-77;
sine[17284]=-77;
sine[17285]=-77;
sine[17286]=-77;
sine[17287]=-77;
sine[17288]=-77;
sine[17289]=-77;
sine[17290]=-77;
sine[17291]=-77;
sine[17292]=-77;
sine[17293]=-77;
sine[17294]=-77;
sine[17295]=-77;
sine[17296]=-77;
sine[17297]=-77;
sine[17298]=-77;
sine[17299]=-78;
sine[17300]=-78;
sine[17301]=-78;
sine[17302]=-78;
sine[17303]=-78;
sine[17304]=-78;
sine[17305]=-78;
sine[17306]=-78;
sine[17307]=-78;
sine[17308]=-78;
sine[17309]=-78;
sine[17310]=-78;
sine[17311]=-78;
sine[17312]=-78;
sine[17313]=-78;
sine[17314]=-78;
sine[17315]=-78;
sine[17316]=-78;
sine[17317]=-78;
sine[17318]=-78;
sine[17319]=-78;
sine[17320]=-78;
sine[17321]=-78;
sine[17322]=-78;
sine[17323]=-78;
sine[17324]=-78;
sine[17325]=-78;
sine[17326]=-78;
sine[17327]=-78;
sine[17328]=-78;
sine[17329]=-78;
sine[17330]=-78;
sine[17331]=-78;
sine[17332]=-78;
sine[17333]=-78;
sine[17334]=-78;
sine[17335]=-78;
sine[17336]=-78;
sine[17337]=-78;
sine[17338]=-78;
sine[17339]=-78;
sine[17340]=-78;
sine[17341]=-78;
sine[17342]=-78;
sine[17343]=-78;
sine[17344]=-78;
sine[17345]=-78;
sine[17346]=-78;
sine[17347]=-78;
sine[17348]=-78;
sine[17349]=-78;
sine[17350]=-78;
sine[17351]=-78;
sine[17352]=-78;
sine[17353]=-78;
sine[17354]=-78;
sine[17355]=-78;
sine[17356]=-78;
sine[17357]=-78;
sine[17358]=-78;
sine[17359]=-78;
sine[17360]=-78;
sine[17361]=-78;
sine[17362]=-78;
sine[17363]=-78;
sine[17364]=-78;
sine[17365]=-78;
sine[17366]=-78;
sine[17367]=-78;
sine[17368]=-78;
sine[17369]=-78;
sine[17370]=-78;
sine[17371]=-78;
sine[17372]=-78;
sine[17373]=-78;
sine[17374]=-78;
sine[17375]=-78;
sine[17376]=-78;
sine[17377]=-78;
sine[17378]=-78;
sine[17379]=-78;
sine[17380]=-78;
sine[17381]=-78;
sine[17382]=-78;
sine[17383]=-78;
sine[17384]=-78;
sine[17385]=-78;
sine[17386]=-78;
sine[17387]=-78;
sine[17388]=-78;
sine[17389]=-78;
sine[17390]=-78;
sine[17391]=-78;
sine[17392]=-78;
sine[17393]=-78;
sine[17394]=-78;
sine[17395]=-78;
sine[17396]=-78;
sine[17397]=-78;
sine[17398]=-78;
sine[17399]=-78;
sine[17400]=-78;
sine[17401]=-78;
sine[17402]=-78;
sine[17403]=-78;
sine[17404]=-78;
sine[17405]=-78;
sine[17406]=-78;
sine[17407]=-78;
sine[17408]=-78;
sine[17409]=-78;
sine[17410]=-78;
sine[17411]=-78;
sine[17412]=-78;
sine[17413]=-78;
sine[17414]=-78;
sine[17415]=-78;
sine[17416]=-78;
sine[17417]=-78;
sine[17418]=-78;
sine[17419]=-78;
sine[17420]=-78;
sine[17421]=-78;
sine[17422]=-78;
sine[17423]=-78;
sine[17424]=-78;
sine[17425]=-78;
sine[17426]=-78;
sine[17427]=-78;
sine[17428]=-78;
sine[17429]=-78;
sine[17430]=-78;
sine[17431]=-78;
sine[17432]=-78;
sine[17433]=-78;
sine[17434]=-78;
sine[17435]=-78;
sine[17436]=-78;
sine[17437]=-78;
sine[17438]=-78;
sine[17439]=-78;
sine[17440]=-78;
sine[17441]=-78;
sine[17442]=-78;
sine[17443]=-78;
sine[17444]=-78;
sine[17445]=-78;
sine[17446]=-78;
sine[17447]=-78;
sine[17448]=-78;
sine[17449]=-78;
sine[17450]=-78;
sine[17451]=-78;
sine[17452]=-78;
sine[17453]=-78;
sine[17454]=-78;
sine[17455]=-78;
sine[17456]=-78;
sine[17457]=-78;
sine[17458]=-78;
sine[17459]=-78;
sine[17460]=-78;
sine[17461]=-78;
sine[17462]=-78;
sine[17463]=-78;
sine[17464]=-78;
sine[17465]=-78;
sine[17466]=-78;
sine[17467]=-78;
sine[17468]=-78;
sine[17469]=-78;
sine[17470]=-78;
sine[17471]=-78;
sine[17472]=-78;
sine[17473]=-78;
sine[17474]=-78;
sine[17475]=-78;
sine[17476]=-78;
sine[17477]=-78;
sine[17478]=-78;
sine[17479]=-78;
sine[17480]=-78;
sine[17481]=-78;
sine[17482]=-78;
sine[17483]=-78;
sine[17484]=-78;
sine[17485]=-78;
sine[17486]=-78;
sine[17487]=-78;
sine[17488]=-78;
sine[17489]=-78;
sine[17490]=-78;
sine[17491]=-78;
sine[17492]=-78;
sine[17493]=-78;
sine[17494]=-78;
sine[17495]=-78;
sine[17496]=-78;
sine[17497]=-78;
sine[17498]=-78;
sine[17499]=-78;
sine[17500]=-78;
sine[17501]=-78;
sine[17502]=-78;
sine[17503]=-78;
sine[17504]=-78;
sine[17505]=-78;
sine[17506]=-78;
sine[17507]=-78;
sine[17508]=-78;
sine[17509]=-78;
sine[17510]=-78;
sine[17511]=-78;
sine[17512]=-78;
sine[17513]=-78;
sine[17514]=-78;
sine[17515]=-78;
sine[17516]=-78;
sine[17517]=-78;
sine[17518]=-78;
sine[17519]=-78;
sine[17520]=-78;
sine[17521]=-78;
sine[17522]=-78;
sine[17523]=-78;
sine[17524]=-78;
sine[17525]=-78;
sine[17526]=-78;
sine[17527]=-78;
sine[17528]=-78;
sine[17529]=-78;
sine[17530]=-78;
sine[17531]=-78;
sine[17532]=-78;
sine[17533]=-78;
sine[17534]=-78;
sine[17535]=-78;
sine[17536]=-78;
sine[17537]=-78;
sine[17538]=-78;
sine[17539]=-78;
sine[17540]=-78;
sine[17541]=-78;
sine[17542]=-78;
sine[17543]=-78;
sine[17544]=-78;
sine[17545]=-78;
sine[17546]=-78;
sine[17547]=-78;
sine[17548]=-78;
sine[17549]=-78;
sine[17550]=-78;
sine[17551]=-78;
sine[17552]=-78;
sine[17553]=-78;
sine[17554]=-78;
sine[17555]=-78;
sine[17556]=-78;
sine[17557]=-78;
sine[17558]=-78;
sine[17559]=-78;
sine[17560]=-78;
sine[17561]=-78;
sine[17562]=-78;
sine[17563]=-78;
sine[17564]=-78;
sine[17565]=-78;
sine[17566]=-78;
sine[17567]=-78;
sine[17568]=-78;
sine[17569]=-78;
sine[17570]=-78;
sine[17571]=-78;
sine[17572]=-78;
sine[17573]=-78;
sine[17574]=-78;
sine[17575]=-78;
sine[17576]=-78;
sine[17577]=-78;
sine[17578]=-78;
sine[17579]=-78;
sine[17580]=-78;
sine[17581]=-78;
sine[17582]=-78;
sine[17583]=-78;
sine[17584]=-78;
sine[17585]=-78;
sine[17586]=-78;
sine[17587]=-78;
sine[17588]=-78;
sine[17589]=-78;
sine[17590]=-78;
sine[17591]=-78;
sine[17592]=-78;
sine[17593]=-78;
sine[17594]=-78;
sine[17595]=-78;
sine[17596]=-78;
sine[17597]=-78;
sine[17598]=-78;
sine[17599]=-78;
sine[17600]=-78;
sine[17601]=-78;
sine[17602]=-78;
sine[17603]=-78;
sine[17604]=-78;
sine[17605]=-78;
sine[17606]=-78;
sine[17607]=-78;
sine[17608]=-78;
sine[17609]=-78;
sine[17610]=-78;
sine[17611]=-78;
sine[17612]=-78;
sine[17613]=-78;
sine[17614]=-78;
sine[17615]=-78;
sine[17616]=-78;
sine[17617]=-78;
sine[17618]=-78;
sine[17619]=-78;
sine[17620]=-78;
sine[17621]=-78;
sine[17622]=-78;
sine[17623]=-78;
sine[17624]=-78;
sine[17625]=-78;
sine[17626]=-78;
sine[17627]=-78;
sine[17628]=-78;
sine[17629]=-78;
sine[17630]=-78;
sine[17631]=-78;
sine[17632]=-78;
sine[17633]=-78;
sine[17634]=-78;
sine[17635]=-78;
sine[17636]=-78;
sine[17637]=-78;
sine[17638]=-78;
sine[17639]=-78;
sine[17640]=-78;
sine[17641]=-78;
sine[17642]=-78;
sine[17643]=-78;
sine[17644]=-78;
sine[17645]=-78;
sine[17646]=-78;
sine[17647]=-78;
sine[17648]=-78;
sine[17649]=-78;
sine[17650]=-78;
sine[17651]=-78;
sine[17652]=-78;
sine[17653]=-78;
sine[17654]=-78;
sine[17655]=-78;
sine[17656]=-78;
sine[17657]=-78;
sine[17658]=-78;
sine[17659]=-78;
sine[17660]=-78;
sine[17661]=-78;
sine[17662]=-78;
sine[17663]=-78;
sine[17664]=-78;
sine[17665]=-78;
sine[17666]=-78;
sine[17667]=-78;
sine[17668]=-78;
sine[17669]=-78;
sine[17670]=-78;
sine[17671]=-78;
sine[17672]=-78;
sine[17673]=-78;
sine[17674]=-78;
sine[17675]=-78;
sine[17676]=-78;
sine[17677]=-78;
sine[17678]=-78;
sine[17679]=-78;
sine[17680]=-78;
sine[17681]=-78;
sine[17682]=-78;
sine[17683]=-78;
sine[17684]=-78;
sine[17685]=-78;
sine[17686]=-78;
sine[17687]=-78;
sine[17688]=-78;
sine[17689]=-78;
sine[17690]=-78;
sine[17691]=-78;
sine[17692]=-78;
sine[17693]=-78;
sine[17694]=-78;
sine[17695]=-78;
sine[17696]=-78;
sine[17697]=-78;
sine[17698]=-78;
sine[17699]=-78;
sine[17700]=-78;
sine[17701]=-78;
sine[17702]=-77;
sine[17703]=-77;
sine[17704]=-77;
sine[17705]=-77;
sine[17706]=-77;
sine[17707]=-77;
sine[17708]=-77;
sine[17709]=-77;
sine[17710]=-77;
sine[17711]=-77;
sine[17712]=-77;
sine[17713]=-77;
sine[17714]=-77;
sine[17715]=-77;
sine[17716]=-77;
sine[17717]=-77;
sine[17718]=-77;
sine[17719]=-77;
sine[17720]=-77;
sine[17721]=-77;
sine[17722]=-77;
sine[17723]=-77;
sine[17724]=-77;
sine[17725]=-77;
sine[17726]=-77;
sine[17727]=-77;
sine[17728]=-77;
sine[17729]=-77;
sine[17730]=-77;
sine[17731]=-77;
sine[17732]=-77;
sine[17733]=-77;
sine[17734]=-77;
sine[17735]=-77;
sine[17736]=-77;
sine[17737]=-77;
sine[17738]=-77;
sine[17739]=-77;
sine[17740]=-77;
sine[17741]=-77;
sine[17742]=-77;
sine[17743]=-77;
sine[17744]=-77;
sine[17745]=-77;
sine[17746]=-77;
sine[17747]=-77;
sine[17748]=-77;
sine[17749]=-77;
sine[17750]=-77;
sine[17751]=-77;
sine[17752]=-77;
sine[17753]=-77;
sine[17754]=-77;
sine[17755]=-77;
sine[17756]=-77;
sine[17757]=-77;
sine[17758]=-77;
sine[17759]=-77;
sine[17760]=-77;
sine[17761]=-77;
sine[17762]=-77;
sine[17763]=-77;
sine[17764]=-77;
sine[17765]=-77;
sine[17766]=-77;
sine[17767]=-77;
sine[17768]=-77;
sine[17769]=-77;
sine[17770]=-77;
sine[17771]=-77;
sine[17772]=-77;
sine[17773]=-77;
sine[17774]=-77;
sine[17775]=-77;
sine[17776]=-77;
sine[17777]=-77;
sine[17778]=-77;
sine[17779]=-77;
sine[17780]=-77;
sine[17781]=-77;
sine[17782]=-77;
sine[17783]=-77;
sine[17784]=-77;
sine[17785]=-77;
sine[17786]=-77;
sine[17787]=-77;
sine[17788]=-77;
sine[17789]=-77;
sine[17790]=-77;
sine[17791]=-77;
sine[17792]=-77;
sine[17793]=-77;
sine[17794]=-77;
sine[17795]=-77;
sine[17796]=-77;
sine[17797]=-77;
sine[17798]=-77;
sine[17799]=-77;
sine[17800]=-77;
sine[17801]=-77;
sine[17802]=-77;
sine[17803]=-77;
sine[17804]=-77;
sine[17805]=-77;
sine[17806]=-77;
sine[17807]=-77;
sine[17808]=-77;
sine[17809]=-77;
sine[17810]=-77;
sine[17811]=-77;
sine[17812]=-77;
sine[17813]=-77;
sine[17814]=-77;
sine[17815]=-77;
sine[17816]=-77;
sine[17817]=-77;
sine[17818]=-77;
sine[17819]=-77;
sine[17820]=-77;
sine[17821]=-77;
sine[17822]=-77;
sine[17823]=-77;
sine[17824]=-77;
sine[17825]=-77;
sine[17826]=-76;
sine[17827]=-76;
sine[17828]=-76;
sine[17829]=-76;
sine[17830]=-76;
sine[17831]=-76;
sine[17832]=-76;
sine[17833]=-76;
sine[17834]=-76;
sine[17835]=-76;
sine[17836]=-76;
sine[17837]=-76;
sine[17838]=-76;
sine[17839]=-76;
sine[17840]=-76;
sine[17841]=-76;
sine[17842]=-76;
sine[17843]=-76;
sine[17844]=-76;
sine[17845]=-76;
sine[17846]=-76;
sine[17847]=-76;
sine[17848]=-76;
sine[17849]=-76;
sine[17850]=-76;
sine[17851]=-76;
sine[17852]=-76;
sine[17853]=-76;
sine[17854]=-76;
sine[17855]=-76;
sine[17856]=-76;
sine[17857]=-76;
sine[17858]=-76;
sine[17859]=-76;
sine[17860]=-76;
sine[17861]=-76;
sine[17862]=-76;
sine[17863]=-76;
sine[17864]=-76;
sine[17865]=-76;
sine[17866]=-76;
sine[17867]=-76;
sine[17868]=-76;
sine[17869]=-76;
sine[17870]=-76;
sine[17871]=-76;
sine[17872]=-76;
sine[17873]=-76;
sine[17874]=-76;
sine[17875]=-76;
sine[17876]=-76;
sine[17877]=-76;
sine[17878]=-76;
sine[17879]=-76;
sine[17880]=-76;
sine[17881]=-76;
sine[17882]=-76;
sine[17883]=-76;
sine[17884]=-76;
sine[17885]=-76;
sine[17886]=-76;
sine[17887]=-76;
sine[17888]=-76;
sine[17889]=-76;
sine[17890]=-76;
sine[17891]=-76;
sine[17892]=-76;
sine[17893]=-76;
sine[17894]=-76;
sine[17895]=-76;
sine[17896]=-76;
sine[17897]=-76;
sine[17898]=-76;
sine[17899]=-76;
sine[17900]=-76;
sine[17901]=-76;
sine[17902]=-76;
sine[17903]=-76;
sine[17904]=-76;
sine[17905]=-76;
sine[17906]=-76;
sine[17907]=-76;
sine[17908]=-76;
sine[17909]=-76;
sine[17910]=-76;
sine[17911]=-76;
sine[17912]=-76;
sine[17913]=-76;
sine[17914]=-75;
sine[17915]=-75;
sine[17916]=-75;
sine[17917]=-75;
sine[17918]=-75;
sine[17919]=-75;
sine[17920]=-75;
sine[17921]=-75;
sine[17922]=-75;
sine[17923]=-75;
sine[17924]=-75;
sine[17925]=-75;
sine[17926]=-75;
sine[17927]=-75;
sine[17928]=-75;
sine[17929]=-75;
sine[17930]=-75;
sine[17931]=-75;
sine[17932]=-75;
sine[17933]=-75;
sine[17934]=-75;
sine[17935]=-75;
sine[17936]=-75;
sine[17937]=-75;
sine[17938]=-75;
sine[17939]=-75;
sine[17940]=-75;
sine[17941]=-75;
sine[17942]=-75;
sine[17943]=-75;
sine[17944]=-75;
sine[17945]=-75;
sine[17946]=-75;
sine[17947]=-75;
sine[17948]=-75;
sine[17949]=-75;
sine[17950]=-75;
sine[17951]=-75;
sine[17952]=-75;
sine[17953]=-75;
sine[17954]=-75;
sine[17955]=-75;
sine[17956]=-75;
sine[17957]=-75;
sine[17958]=-75;
sine[17959]=-75;
sine[17960]=-75;
sine[17961]=-75;
sine[17962]=-75;
sine[17963]=-75;
sine[17964]=-75;
sine[17965]=-75;
sine[17966]=-75;
sine[17967]=-75;
sine[17968]=-75;
sine[17969]=-75;
sine[17970]=-75;
sine[17971]=-75;
sine[17972]=-75;
sine[17973]=-75;
sine[17974]=-75;
sine[17975]=-75;
sine[17976]=-75;
sine[17977]=-75;
sine[17978]=-75;
sine[17979]=-75;
sine[17980]=-75;
sine[17981]=-75;
sine[17982]=-75;
sine[17983]=-75;
sine[17984]=-75;
sine[17985]=-75;
sine[17986]=-75;
sine[17987]=-74;
sine[17988]=-74;
sine[17989]=-74;
sine[17990]=-74;
sine[17991]=-74;
sine[17992]=-74;
sine[17993]=-74;
sine[17994]=-74;
sine[17995]=-74;
sine[17996]=-74;
sine[17997]=-74;
sine[17998]=-74;
sine[17999]=-74;
sine[18000]=-74;
sine[18001]=-74;
sine[18002]=-74;
sine[18003]=-74;
sine[18004]=-74;
sine[18005]=-74;
sine[18006]=-74;
sine[18007]=-74;
sine[18008]=-74;
sine[18009]=-74;
sine[18010]=-74;
sine[18011]=-74;
sine[18012]=-74;
sine[18013]=-74;
sine[18014]=-74;
sine[18015]=-74;
sine[18016]=-74;
sine[18017]=-74;
sine[18018]=-74;
sine[18019]=-74;
sine[18020]=-74;
sine[18021]=-74;
sine[18022]=-74;
sine[18023]=-74;
sine[18024]=-74;
sine[18025]=-74;
sine[18026]=-74;
sine[18027]=-74;
sine[18028]=-74;
sine[18029]=-74;
sine[18030]=-74;
sine[18031]=-74;
sine[18032]=-74;
sine[18033]=-74;
sine[18034]=-74;
sine[18035]=-74;
sine[18036]=-74;
sine[18037]=-74;
sine[18038]=-74;
sine[18039]=-74;
sine[18040]=-74;
sine[18041]=-74;
sine[18042]=-74;
sine[18043]=-74;
sine[18044]=-74;
sine[18045]=-74;
sine[18046]=-74;
sine[18047]=-74;
sine[18048]=-74;
sine[18049]=-74;
sine[18050]=-74;
sine[18051]=-73;
sine[18052]=-73;
sine[18053]=-73;
sine[18054]=-73;
sine[18055]=-73;
sine[18056]=-73;
sine[18057]=-73;
sine[18058]=-73;
sine[18059]=-73;
sine[18060]=-73;
sine[18061]=-73;
sine[18062]=-73;
sine[18063]=-73;
sine[18064]=-73;
sine[18065]=-73;
sine[18066]=-73;
sine[18067]=-73;
sine[18068]=-73;
sine[18069]=-73;
sine[18070]=-73;
sine[18071]=-73;
sine[18072]=-73;
sine[18073]=-73;
sine[18074]=-73;
sine[18075]=-73;
sine[18076]=-73;
sine[18077]=-73;
sine[18078]=-73;
sine[18079]=-73;
sine[18080]=-73;
sine[18081]=-73;
sine[18082]=-73;
sine[18083]=-73;
sine[18084]=-73;
sine[18085]=-73;
sine[18086]=-73;
sine[18087]=-73;
sine[18088]=-73;
sine[18089]=-73;
sine[18090]=-73;
sine[18091]=-73;
sine[18092]=-73;
sine[18093]=-73;
sine[18094]=-73;
sine[18095]=-73;
sine[18096]=-73;
sine[18097]=-73;
sine[18098]=-73;
sine[18099]=-73;
sine[18100]=-73;
sine[18101]=-73;
sine[18102]=-73;
sine[18103]=-73;
sine[18104]=-73;
sine[18105]=-73;
sine[18106]=-73;
sine[18107]=-73;
sine[18108]=-72;
sine[18109]=-72;
sine[18110]=-72;
sine[18111]=-72;
sine[18112]=-72;
sine[18113]=-72;
sine[18114]=-72;
sine[18115]=-72;
sine[18116]=-72;
sine[18117]=-72;
sine[18118]=-72;
sine[18119]=-72;
sine[18120]=-72;
sine[18121]=-72;
sine[18122]=-72;
sine[18123]=-72;
sine[18124]=-72;
sine[18125]=-72;
sine[18126]=-72;
sine[18127]=-72;
sine[18128]=-72;
sine[18129]=-72;
sine[18130]=-72;
sine[18131]=-72;
sine[18132]=-72;
sine[18133]=-72;
sine[18134]=-72;
sine[18135]=-72;
sine[18136]=-72;
sine[18137]=-72;
sine[18138]=-72;
sine[18139]=-72;
sine[18140]=-72;
sine[18141]=-72;
sine[18142]=-72;
sine[18143]=-72;
sine[18144]=-72;
sine[18145]=-72;
sine[18146]=-72;
sine[18147]=-72;
sine[18148]=-72;
sine[18149]=-72;
sine[18150]=-72;
sine[18151]=-72;
sine[18152]=-72;
sine[18153]=-72;
sine[18154]=-72;
sine[18155]=-72;
sine[18156]=-72;
sine[18157]=-72;
sine[18158]=-72;
sine[18159]=-72;
sine[18160]=-72;
sine[18161]=-71;
sine[18162]=-71;
sine[18163]=-71;
sine[18164]=-71;
sine[18165]=-71;
sine[18166]=-71;
sine[18167]=-71;
sine[18168]=-71;
sine[18169]=-71;
sine[18170]=-71;
sine[18171]=-71;
sine[18172]=-71;
sine[18173]=-71;
sine[18174]=-71;
sine[18175]=-71;
sine[18176]=-71;
sine[18177]=-71;
sine[18178]=-71;
sine[18179]=-71;
sine[18180]=-71;
sine[18181]=-71;
sine[18182]=-71;
sine[18183]=-71;
sine[18184]=-71;
sine[18185]=-71;
sine[18186]=-71;
sine[18187]=-71;
sine[18188]=-71;
sine[18189]=-71;
sine[18190]=-71;
sine[18191]=-71;
sine[18192]=-71;
sine[18193]=-71;
sine[18194]=-71;
sine[18195]=-71;
sine[18196]=-71;
sine[18197]=-71;
sine[18198]=-71;
sine[18199]=-71;
sine[18200]=-71;
sine[18201]=-71;
sine[18202]=-71;
sine[18203]=-71;
sine[18204]=-71;
sine[18205]=-71;
sine[18206]=-71;
sine[18207]=-71;
sine[18208]=-71;
sine[18209]=-71;
sine[18210]=-70;
sine[18211]=-70;
sine[18212]=-70;
sine[18213]=-70;
sine[18214]=-70;
sine[18215]=-70;
sine[18216]=-70;
sine[18217]=-70;
sine[18218]=-70;
sine[18219]=-70;
sine[18220]=-70;
sine[18221]=-70;
sine[18222]=-70;
sine[18223]=-70;
sine[18224]=-70;
sine[18225]=-70;
sine[18226]=-70;
sine[18227]=-70;
sine[18228]=-70;
sine[18229]=-70;
sine[18230]=-70;
sine[18231]=-70;
sine[18232]=-70;
sine[18233]=-70;
sine[18234]=-70;
sine[18235]=-70;
sine[18236]=-70;
sine[18237]=-70;
sine[18238]=-70;
sine[18239]=-70;
sine[18240]=-70;
sine[18241]=-70;
sine[18242]=-70;
sine[18243]=-70;
sine[18244]=-70;
sine[18245]=-70;
sine[18246]=-70;
sine[18247]=-70;
sine[18248]=-70;
sine[18249]=-70;
sine[18250]=-70;
sine[18251]=-70;
sine[18252]=-70;
sine[18253]=-70;
sine[18254]=-70;
sine[18255]=-69;
sine[18256]=-69;
sine[18257]=-69;
sine[18258]=-69;
sine[18259]=-69;
sine[18260]=-69;
sine[18261]=-69;
sine[18262]=-69;
sine[18263]=-69;
sine[18264]=-69;
sine[18265]=-69;
sine[18266]=-69;
sine[18267]=-69;
sine[18268]=-69;
sine[18269]=-69;
sine[18270]=-69;
sine[18271]=-69;
sine[18272]=-69;
sine[18273]=-69;
sine[18274]=-69;
sine[18275]=-69;
sine[18276]=-69;
sine[18277]=-69;
sine[18278]=-69;
sine[18279]=-69;
sine[18280]=-69;
sine[18281]=-69;
sine[18282]=-69;
sine[18283]=-69;
sine[18284]=-69;
sine[18285]=-69;
sine[18286]=-69;
sine[18287]=-69;
sine[18288]=-69;
sine[18289]=-69;
sine[18290]=-69;
sine[18291]=-69;
sine[18292]=-69;
sine[18293]=-69;
sine[18294]=-69;
sine[18295]=-69;
sine[18296]=-69;
sine[18297]=-69;
sine[18298]=-69;
sine[18299]=-68;
sine[18300]=-68;
sine[18301]=-68;
sine[18302]=-68;
sine[18303]=-68;
sine[18304]=-68;
sine[18305]=-68;
sine[18306]=-68;
sine[18307]=-68;
sine[18308]=-68;
sine[18309]=-68;
sine[18310]=-68;
sine[18311]=-68;
sine[18312]=-68;
sine[18313]=-68;
sine[18314]=-68;
sine[18315]=-68;
sine[18316]=-68;
sine[18317]=-68;
sine[18318]=-68;
sine[18319]=-68;
sine[18320]=-68;
sine[18321]=-68;
sine[18322]=-68;
sine[18323]=-68;
sine[18324]=-68;
sine[18325]=-68;
sine[18326]=-68;
sine[18327]=-68;
sine[18328]=-68;
sine[18329]=-68;
sine[18330]=-68;
sine[18331]=-68;
sine[18332]=-68;
sine[18333]=-68;
sine[18334]=-68;
sine[18335]=-68;
sine[18336]=-68;
sine[18337]=-68;
sine[18338]=-68;
sine[18339]=-68;
sine[18340]=-67;
sine[18341]=-67;
sine[18342]=-67;
sine[18343]=-67;
sine[18344]=-67;
sine[18345]=-67;
sine[18346]=-67;
sine[18347]=-67;
sine[18348]=-67;
sine[18349]=-67;
sine[18350]=-67;
sine[18351]=-67;
sine[18352]=-67;
sine[18353]=-67;
sine[18354]=-67;
sine[18355]=-67;
sine[18356]=-67;
sine[18357]=-67;
sine[18358]=-67;
sine[18359]=-67;
sine[18360]=-67;
sine[18361]=-67;
sine[18362]=-67;
sine[18363]=-67;
sine[18364]=-67;
sine[18365]=-67;
sine[18366]=-67;
sine[18367]=-67;
sine[18368]=-67;
sine[18369]=-67;
sine[18370]=-67;
sine[18371]=-67;
sine[18372]=-67;
sine[18373]=-67;
sine[18374]=-67;
sine[18375]=-67;
sine[18376]=-67;
sine[18377]=-67;
sine[18378]=-67;
sine[18379]=-67;
sine[18380]=-66;
sine[18381]=-66;
sine[18382]=-66;
sine[18383]=-66;
sine[18384]=-66;
sine[18385]=-66;
sine[18386]=-66;
sine[18387]=-66;
sine[18388]=-66;
sine[18389]=-66;
sine[18390]=-66;
sine[18391]=-66;
sine[18392]=-66;
sine[18393]=-66;
sine[18394]=-66;
sine[18395]=-66;
sine[18396]=-66;
sine[18397]=-66;
sine[18398]=-66;
sine[18399]=-66;
sine[18400]=-66;
sine[18401]=-66;
sine[18402]=-66;
sine[18403]=-66;
sine[18404]=-66;
sine[18405]=-66;
sine[18406]=-66;
sine[18407]=-66;
sine[18408]=-66;
sine[18409]=-66;
sine[18410]=-66;
sine[18411]=-66;
sine[18412]=-66;
sine[18413]=-66;
sine[18414]=-66;
sine[18415]=-66;
sine[18416]=-66;
sine[18417]=-66;
sine[18418]=-65;
sine[18419]=-65;
sine[18420]=-65;
sine[18421]=-65;
sine[18422]=-65;
sine[18423]=-65;
sine[18424]=-65;
sine[18425]=-65;
sine[18426]=-65;
sine[18427]=-65;
sine[18428]=-65;
sine[18429]=-65;
sine[18430]=-65;
sine[18431]=-65;
sine[18432]=-65;
sine[18433]=-65;
sine[18434]=-65;
sine[18435]=-65;
sine[18436]=-65;
sine[18437]=-65;
sine[18438]=-65;
sine[18439]=-65;
sine[18440]=-65;
sine[18441]=-65;
sine[18442]=-65;
sine[18443]=-65;
sine[18444]=-65;
sine[18445]=-65;
sine[18446]=-65;
sine[18447]=-65;
sine[18448]=-65;
sine[18449]=-65;
sine[18450]=-65;
sine[18451]=-65;
sine[18452]=-65;
sine[18453]=-65;
sine[18454]=-65;
sine[18455]=-64;
sine[18456]=-64;
sine[18457]=-64;
sine[18458]=-64;
sine[18459]=-64;
sine[18460]=-64;
sine[18461]=-64;
sine[18462]=-64;
sine[18463]=-64;
sine[18464]=-64;
sine[18465]=-64;
sine[18466]=-64;
sine[18467]=-64;
sine[18468]=-64;
sine[18469]=-64;
sine[18470]=-64;
sine[18471]=-64;
sine[18472]=-64;
sine[18473]=-64;
sine[18474]=-64;
sine[18475]=-64;
sine[18476]=-64;
sine[18477]=-64;
sine[18478]=-64;
sine[18479]=-64;
sine[18480]=-64;
sine[18481]=-64;
sine[18482]=-64;
sine[18483]=-64;
sine[18484]=-64;
sine[18485]=-64;
sine[18486]=-64;
sine[18487]=-64;
sine[18488]=-64;
sine[18489]=-64;
sine[18490]=-63;
sine[18491]=-63;
sine[18492]=-63;
sine[18493]=-63;
sine[18494]=-63;
sine[18495]=-63;
sine[18496]=-63;
sine[18497]=-63;
sine[18498]=-63;
sine[18499]=-63;
sine[18500]=-63;
sine[18501]=-63;
sine[18502]=-63;
sine[18503]=-63;
sine[18504]=-63;
sine[18505]=-63;
sine[18506]=-63;
sine[18507]=-63;
sine[18508]=-63;
sine[18509]=-63;
sine[18510]=-63;
sine[18511]=-63;
sine[18512]=-63;
sine[18513]=-63;
sine[18514]=-63;
sine[18515]=-63;
sine[18516]=-63;
sine[18517]=-63;
sine[18518]=-63;
sine[18519]=-63;
sine[18520]=-63;
sine[18521]=-63;
sine[18522]=-63;
sine[18523]=-63;
sine[18524]=-63;
sine[18525]=-62;
sine[18526]=-62;
sine[18527]=-62;
sine[18528]=-62;
sine[18529]=-62;
sine[18530]=-62;
sine[18531]=-62;
sine[18532]=-62;
sine[18533]=-62;
sine[18534]=-62;
sine[18535]=-62;
sine[18536]=-62;
sine[18537]=-62;
sine[18538]=-62;
sine[18539]=-62;
sine[18540]=-62;
sine[18541]=-62;
sine[18542]=-62;
sine[18543]=-62;
sine[18544]=-62;
sine[18545]=-62;
sine[18546]=-62;
sine[18547]=-62;
sine[18548]=-62;
sine[18549]=-62;
sine[18550]=-62;
sine[18551]=-62;
sine[18552]=-62;
sine[18553]=-62;
sine[18554]=-62;
sine[18555]=-62;
sine[18556]=-62;
sine[18557]=-62;
sine[18558]=-61;
sine[18559]=-61;
sine[18560]=-61;
sine[18561]=-61;
sine[18562]=-61;
sine[18563]=-61;
sine[18564]=-61;
sine[18565]=-61;
sine[18566]=-61;
sine[18567]=-61;
sine[18568]=-61;
sine[18569]=-61;
sine[18570]=-61;
sine[18571]=-61;
sine[18572]=-61;
sine[18573]=-61;
sine[18574]=-61;
sine[18575]=-61;
sine[18576]=-61;
sine[18577]=-61;
sine[18578]=-61;
sine[18579]=-61;
sine[18580]=-61;
sine[18581]=-61;
sine[18582]=-61;
sine[18583]=-61;
sine[18584]=-61;
sine[18585]=-61;
sine[18586]=-61;
sine[18587]=-61;
sine[18588]=-61;
sine[18589]=-61;
sine[18590]=-61;
sine[18591]=-60;
sine[18592]=-60;
sine[18593]=-60;
sine[18594]=-60;
sine[18595]=-60;
sine[18596]=-60;
sine[18597]=-60;
sine[18598]=-60;
sine[18599]=-60;
sine[18600]=-60;
sine[18601]=-60;
sine[18602]=-60;
sine[18603]=-60;
sine[18604]=-60;
sine[18605]=-60;
sine[18606]=-60;
sine[18607]=-60;
sine[18608]=-60;
sine[18609]=-60;
sine[18610]=-60;
sine[18611]=-60;
sine[18612]=-60;
sine[18613]=-60;
sine[18614]=-60;
sine[18615]=-60;
sine[18616]=-60;
sine[18617]=-60;
sine[18618]=-60;
sine[18619]=-60;
sine[18620]=-60;
sine[18621]=-60;
sine[18622]=-60;
sine[18623]=-59;
sine[18624]=-59;
sine[18625]=-59;
sine[18626]=-59;
sine[18627]=-59;
sine[18628]=-59;
sine[18629]=-59;
sine[18630]=-59;
sine[18631]=-59;
sine[18632]=-59;
sine[18633]=-59;
sine[18634]=-59;
sine[18635]=-59;
sine[18636]=-59;
sine[18637]=-59;
sine[18638]=-59;
sine[18639]=-59;
sine[18640]=-59;
sine[18641]=-59;
sine[18642]=-59;
sine[18643]=-59;
sine[18644]=-59;
sine[18645]=-59;
sine[18646]=-59;
sine[18647]=-59;
sine[18648]=-59;
sine[18649]=-59;
sine[18650]=-59;
sine[18651]=-59;
sine[18652]=-59;
sine[18653]=-59;
sine[18654]=-58;
sine[18655]=-58;
sine[18656]=-58;
sine[18657]=-58;
sine[18658]=-58;
sine[18659]=-58;
sine[18660]=-58;
sine[18661]=-58;
sine[18662]=-58;
sine[18663]=-58;
sine[18664]=-58;
sine[18665]=-58;
sine[18666]=-58;
sine[18667]=-58;
sine[18668]=-58;
sine[18669]=-58;
sine[18670]=-58;
sine[18671]=-58;
sine[18672]=-58;
sine[18673]=-58;
sine[18674]=-58;
sine[18675]=-58;
sine[18676]=-58;
sine[18677]=-58;
sine[18678]=-58;
sine[18679]=-58;
sine[18680]=-58;
sine[18681]=-58;
sine[18682]=-58;
sine[18683]=-58;
sine[18684]=-57;
sine[18685]=-57;
sine[18686]=-57;
sine[18687]=-57;
sine[18688]=-57;
sine[18689]=-57;
sine[18690]=-57;
sine[18691]=-57;
sine[18692]=-57;
sine[18693]=-57;
sine[18694]=-57;
sine[18695]=-57;
sine[18696]=-57;
sine[18697]=-57;
sine[18698]=-57;
sine[18699]=-57;
sine[18700]=-57;
sine[18701]=-57;
sine[18702]=-57;
sine[18703]=-57;
sine[18704]=-57;
sine[18705]=-57;
sine[18706]=-57;
sine[18707]=-57;
sine[18708]=-57;
sine[18709]=-57;
sine[18710]=-57;
sine[18711]=-57;
sine[18712]=-57;
sine[18713]=-57;
sine[18714]=-56;
sine[18715]=-56;
sine[18716]=-56;
sine[18717]=-56;
sine[18718]=-56;
sine[18719]=-56;
sine[18720]=-56;
sine[18721]=-56;
sine[18722]=-56;
sine[18723]=-56;
sine[18724]=-56;
sine[18725]=-56;
sine[18726]=-56;
sine[18727]=-56;
sine[18728]=-56;
sine[18729]=-56;
sine[18730]=-56;
sine[18731]=-56;
sine[18732]=-56;
sine[18733]=-56;
sine[18734]=-56;
sine[18735]=-56;
sine[18736]=-56;
sine[18737]=-56;
sine[18738]=-56;
sine[18739]=-56;
sine[18740]=-56;
sine[18741]=-56;
sine[18742]=-56;
sine[18743]=-55;
sine[18744]=-55;
sine[18745]=-55;
sine[18746]=-55;
sine[18747]=-55;
sine[18748]=-55;
sine[18749]=-55;
sine[18750]=-55;
sine[18751]=-55;
sine[18752]=-55;
sine[18753]=-55;
sine[18754]=-55;
sine[18755]=-55;
sine[18756]=-55;
sine[18757]=-55;
sine[18758]=-55;
sine[18759]=-55;
sine[18760]=-55;
sine[18761]=-55;
sine[18762]=-55;
sine[18763]=-55;
sine[18764]=-55;
sine[18765]=-55;
sine[18766]=-55;
sine[18767]=-55;
sine[18768]=-55;
sine[18769]=-55;
sine[18770]=-55;
sine[18771]=-55;
sine[18772]=-54;
sine[18773]=-54;
sine[18774]=-54;
sine[18775]=-54;
sine[18776]=-54;
sine[18777]=-54;
sine[18778]=-54;
sine[18779]=-54;
sine[18780]=-54;
sine[18781]=-54;
sine[18782]=-54;
sine[18783]=-54;
sine[18784]=-54;
sine[18785]=-54;
sine[18786]=-54;
sine[18787]=-54;
sine[18788]=-54;
sine[18789]=-54;
sine[18790]=-54;
sine[18791]=-54;
sine[18792]=-54;
sine[18793]=-54;
sine[18794]=-54;
sine[18795]=-54;
sine[18796]=-54;
sine[18797]=-54;
sine[18798]=-54;
sine[18799]=-54;
sine[18800]=-53;
sine[18801]=-53;
sine[18802]=-53;
sine[18803]=-53;
sine[18804]=-53;
sine[18805]=-53;
sine[18806]=-53;
sine[18807]=-53;
sine[18808]=-53;
sine[18809]=-53;
sine[18810]=-53;
sine[18811]=-53;
sine[18812]=-53;
sine[18813]=-53;
sine[18814]=-53;
sine[18815]=-53;
sine[18816]=-53;
sine[18817]=-53;
sine[18818]=-53;
sine[18819]=-53;
sine[18820]=-53;
sine[18821]=-53;
sine[18822]=-53;
sine[18823]=-53;
sine[18824]=-53;
sine[18825]=-53;
sine[18826]=-53;
sine[18827]=-53;
sine[18828]=-52;
sine[18829]=-52;
sine[18830]=-52;
sine[18831]=-52;
sine[18832]=-52;
sine[18833]=-52;
sine[18834]=-52;
sine[18835]=-52;
sine[18836]=-52;
sine[18837]=-52;
sine[18838]=-52;
sine[18839]=-52;
sine[18840]=-52;
sine[18841]=-52;
sine[18842]=-52;
sine[18843]=-52;
sine[18844]=-52;
sine[18845]=-52;
sine[18846]=-52;
sine[18847]=-52;
sine[18848]=-52;
sine[18849]=-52;
sine[18850]=-52;
sine[18851]=-52;
sine[18852]=-52;
sine[18853]=-52;
sine[18854]=-52;
sine[18855]=-51;
sine[18856]=-51;
sine[18857]=-51;
sine[18858]=-51;
sine[18859]=-51;
sine[18860]=-51;
sine[18861]=-51;
sine[18862]=-51;
sine[18863]=-51;
sine[18864]=-51;
sine[18865]=-51;
sine[18866]=-51;
sine[18867]=-51;
sine[18868]=-51;
sine[18869]=-51;
sine[18870]=-51;
sine[18871]=-51;
sine[18872]=-51;
sine[18873]=-51;
sine[18874]=-51;
sine[18875]=-51;
sine[18876]=-51;
sine[18877]=-51;
sine[18878]=-51;
sine[18879]=-51;
sine[18880]=-51;
sine[18881]=-51;
sine[18882]=-50;
sine[18883]=-50;
sine[18884]=-50;
sine[18885]=-50;
sine[18886]=-50;
sine[18887]=-50;
sine[18888]=-50;
sine[18889]=-50;
sine[18890]=-50;
sine[18891]=-50;
sine[18892]=-50;
sine[18893]=-50;
sine[18894]=-50;
sine[18895]=-50;
sine[18896]=-50;
sine[18897]=-50;
sine[18898]=-50;
sine[18899]=-50;
sine[18900]=-50;
sine[18901]=-50;
sine[18902]=-50;
sine[18903]=-50;
sine[18904]=-50;
sine[18905]=-50;
sine[18906]=-50;
sine[18907]=-50;
sine[18908]=-49;
sine[18909]=-49;
sine[18910]=-49;
sine[18911]=-49;
sine[18912]=-49;
sine[18913]=-49;
sine[18914]=-49;
sine[18915]=-49;
sine[18916]=-49;
sine[18917]=-49;
sine[18918]=-49;
sine[18919]=-49;
sine[18920]=-49;
sine[18921]=-49;
sine[18922]=-49;
sine[18923]=-49;
sine[18924]=-49;
sine[18925]=-49;
sine[18926]=-49;
sine[18927]=-49;
sine[18928]=-49;
sine[18929]=-49;
sine[18930]=-49;
sine[18931]=-49;
sine[18932]=-49;
sine[18933]=-49;
sine[18934]=-49;
sine[18935]=-48;
sine[18936]=-48;
sine[18937]=-48;
sine[18938]=-48;
sine[18939]=-48;
sine[18940]=-48;
sine[18941]=-48;
sine[18942]=-48;
sine[18943]=-48;
sine[18944]=-48;
sine[18945]=-48;
sine[18946]=-48;
sine[18947]=-48;
sine[18948]=-48;
sine[18949]=-48;
sine[18950]=-48;
sine[18951]=-48;
sine[18952]=-48;
sine[18953]=-48;
sine[18954]=-48;
sine[18955]=-48;
sine[18956]=-48;
sine[18957]=-48;
sine[18958]=-48;
sine[18959]=-48;
sine[18960]=-47;
sine[18961]=-47;
sine[18962]=-47;
sine[18963]=-47;
sine[18964]=-47;
sine[18965]=-47;
sine[18966]=-47;
sine[18967]=-47;
sine[18968]=-47;
sine[18969]=-47;
sine[18970]=-47;
sine[18971]=-47;
sine[18972]=-47;
sine[18973]=-47;
sine[18974]=-47;
sine[18975]=-47;
sine[18976]=-47;
sine[18977]=-47;
sine[18978]=-47;
sine[18979]=-47;
sine[18980]=-47;
sine[18981]=-47;
sine[18982]=-47;
sine[18983]=-47;
sine[18984]=-47;
sine[18985]=-47;
sine[18986]=-46;
sine[18987]=-46;
sine[18988]=-46;
sine[18989]=-46;
sine[18990]=-46;
sine[18991]=-46;
sine[18992]=-46;
sine[18993]=-46;
sine[18994]=-46;
sine[18995]=-46;
sine[18996]=-46;
sine[18997]=-46;
sine[18998]=-46;
sine[18999]=-46;
sine[19000]=-46;
sine[19001]=-46;
sine[19002]=-46;
sine[19003]=-46;
sine[19004]=-46;
sine[19005]=-46;
sine[19006]=-46;
sine[19007]=-46;
sine[19008]=-46;
sine[19009]=-46;
sine[19010]=-46;
sine[19011]=-45;
sine[19012]=-45;
sine[19013]=-45;
sine[19014]=-45;
sine[19015]=-45;
sine[19016]=-45;
sine[19017]=-45;
sine[19018]=-45;
sine[19019]=-45;
sine[19020]=-45;
sine[19021]=-45;
sine[19022]=-45;
sine[19023]=-45;
sine[19024]=-45;
sine[19025]=-45;
sine[19026]=-45;
sine[19027]=-45;
sine[19028]=-45;
sine[19029]=-45;
sine[19030]=-45;
sine[19031]=-45;
sine[19032]=-45;
sine[19033]=-45;
sine[19034]=-45;
sine[19035]=-45;
sine[19036]=-44;
sine[19037]=-44;
sine[19038]=-44;
sine[19039]=-44;
sine[19040]=-44;
sine[19041]=-44;
sine[19042]=-44;
sine[19043]=-44;
sine[19044]=-44;
sine[19045]=-44;
sine[19046]=-44;
sine[19047]=-44;
sine[19048]=-44;
sine[19049]=-44;
sine[19050]=-44;
sine[19051]=-44;
sine[19052]=-44;
sine[19053]=-44;
sine[19054]=-44;
sine[19055]=-44;
sine[19056]=-44;
sine[19057]=-44;
sine[19058]=-44;
sine[19059]=-44;
sine[19060]=-44;
sine[19061]=-43;
sine[19062]=-43;
sine[19063]=-43;
sine[19064]=-43;
sine[19065]=-43;
sine[19066]=-43;
sine[19067]=-43;
sine[19068]=-43;
sine[19069]=-43;
sine[19070]=-43;
sine[19071]=-43;
sine[19072]=-43;
sine[19073]=-43;
sine[19074]=-43;
sine[19075]=-43;
sine[19076]=-43;
sine[19077]=-43;
sine[19078]=-43;
sine[19079]=-43;
sine[19080]=-43;
sine[19081]=-43;
sine[19082]=-43;
sine[19083]=-43;
sine[19084]=-43;
sine[19085]=-42;
sine[19086]=-42;
sine[19087]=-42;
sine[19088]=-42;
sine[19089]=-42;
sine[19090]=-42;
sine[19091]=-42;
sine[19092]=-42;
sine[19093]=-42;
sine[19094]=-42;
sine[19095]=-42;
sine[19096]=-42;
sine[19097]=-42;
sine[19098]=-42;
sine[19099]=-42;
sine[19100]=-42;
sine[19101]=-42;
sine[19102]=-42;
sine[19103]=-42;
sine[19104]=-42;
sine[19105]=-42;
sine[19106]=-42;
sine[19107]=-42;
sine[19108]=-42;
sine[19109]=-41;
sine[19110]=-41;
sine[19111]=-41;
sine[19112]=-41;
sine[19113]=-41;
sine[19114]=-41;
sine[19115]=-41;
sine[19116]=-41;
sine[19117]=-41;
sine[19118]=-41;
sine[19119]=-41;
sine[19120]=-41;
sine[19121]=-41;
sine[19122]=-41;
sine[19123]=-41;
sine[19124]=-41;
sine[19125]=-41;
sine[19126]=-41;
sine[19127]=-41;
sine[19128]=-41;
sine[19129]=-41;
sine[19130]=-41;
sine[19131]=-41;
sine[19132]=-41;
sine[19133]=-40;
sine[19134]=-40;
sine[19135]=-40;
sine[19136]=-40;
sine[19137]=-40;
sine[19138]=-40;
sine[19139]=-40;
sine[19140]=-40;
sine[19141]=-40;
sine[19142]=-40;
sine[19143]=-40;
sine[19144]=-40;
sine[19145]=-40;
sine[19146]=-40;
sine[19147]=-40;
sine[19148]=-40;
sine[19149]=-40;
sine[19150]=-40;
sine[19151]=-40;
sine[19152]=-40;
sine[19153]=-40;
sine[19154]=-40;
sine[19155]=-40;
sine[19156]=-40;
sine[19157]=-39;
sine[19158]=-39;
sine[19159]=-39;
sine[19160]=-39;
sine[19161]=-39;
sine[19162]=-39;
sine[19163]=-39;
sine[19164]=-39;
sine[19165]=-39;
sine[19166]=-39;
sine[19167]=-39;
sine[19168]=-39;
sine[19169]=-39;
sine[19170]=-39;
sine[19171]=-39;
sine[19172]=-39;
sine[19173]=-39;
sine[19174]=-39;
sine[19175]=-39;
sine[19176]=-39;
sine[19177]=-39;
sine[19178]=-39;
sine[19179]=-39;
sine[19180]=-38;
sine[19181]=-38;
sine[19182]=-38;
sine[19183]=-38;
sine[19184]=-38;
sine[19185]=-38;
sine[19186]=-38;
sine[19187]=-38;
sine[19188]=-38;
sine[19189]=-38;
sine[19190]=-38;
sine[19191]=-38;
sine[19192]=-38;
sine[19193]=-38;
sine[19194]=-38;
sine[19195]=-38;
sine[19196]=-38;
sine[19197]=-38;
sine[19198]=-38;
sine[19199]=-38;
sine[19200]=-38;
sine[19201]=-38;
sine[19202]=-38;
sine[19203]=-38;
sine[19204]=-37;
sine[19205]=-37;
sine[19206]=-37;
sine[19207]=-37;
sine[19208]=-37;
sine[19209]=-37;
sine[19210]=-37;
sine[19211]=-37;
sine[19212]=-37;
sine[19213]=-37;
sine[19214]=-37;
sine[19215]=-37;
sine[19216]=-37;
sine[19217]=-37;
sine[19218]=-37;
sine[19219]=-37;
sine[19220]=-37;
sine[19221]=-37;
sine[19222]=-37;
sine[19223]=-37;
sine[19224]=-37;
sine[19225]=-37;
sine[19226]=-37;
sine[19227]=-36;
sine[19228]=-36;
sine[19229]=-36;
sine[19230]=-36;
sine[19231]=-36;
sine[19232]=-36;
sine[19233]=-36;
sine[19234]=-36;
sine[19235]=-36;
sine[19236]=-36;
sine[19237]=-36;
sine[19238]=-36;
sine[19239]=-36;
sine[19240]=-36;
sine[19241]=-36;
sine[19242]=-36;
sine[19243]=-36;
sine[19244]=-36;
sine[19245]=-36;
sine[19246]=-36;
sine[19247]=-36;
sine[19248]=-36;
sine[19249]=-36;
sine[19250]=-35;
sine[19251]=-35;
sine[19252]=-35;
sine[19253]=-35;
sine[19254]=-35;
sine[19255]=-35;
sine[19256]=-35;
sine[19257]=-35;
sine[19258]=-35;
sine[19259]=-35;
sine[19260]=-35;
sine[19261]=-35;
sine[19262]=-35;
sine[19263]=-35;
sine[19264]=-35;
sine[19265]=-35;
sine[19266]=-35;
sine[19267]=-35;
sine[19268]=-35;
sine[19269]=-35;
sine[19270]=-35;
sine[19271]=-35;
sine[19272]=-35;
sine[19273]=-34;
sine[19274]=-34;
sine[19275]=-34;
sine[19276]=-34;
sine[19277]=-34;
sine[19278]=-34;
sine[19279]=-34;
sine[19280]=-34;
sine[19281]=-34;
sine[19282]=-34;
sine[19283]=-34;
sine[19284]=-34;
sine[19285]=-34;
sine[19286]=-34;
sine[19287]=-34;
sine[19288]=-34;
sine[19289]=-34;
sine[19290]=-34;
sine[19291]=-34;
sine[19292]=-34;
sine[19293]=-34;
sine[19294]=-34;
sine[19295]=-33;
sine[19296]=-33;
sine[19297]=-33;
sine[19298]=-33;
sine[19299]=-33;
sine[19300]=-33;
sine[19301]=-33;
sine[19302]=-33;
sine[19303]=-33;
sine[19304]=-33;
sine[19305]=-33;
sine[19306]=-33;
sine[19307]=-33;
sine[19308]=-33;
sine[19309]=-33;
sine[19310]=-33;
sine[19311]=-33;
sine[19312]=-33;
sine[19313]=-33;
sine[19314]=-33;
sine[19315]=-33;
sine[19316]=-33;
sine[19317]=-33;
sine[19318]=-32;
sine[19319]=-32;
sine[19320]=-32;
sine[19321]=-32;
sine[19322]=-32;
sine[19323]=-32;
sine[19324]=-32;
sine[19325]=-32;
sine[19326]=-32;
sine[19327]=-32;
sine[19328]=-32;
sine[19329]=-32;
sine[19330]=-32;
sine[19331]=-32;
sine[19332]=-32;
sine[19333]=-32;
sine[19334]=-32;
sine[19335]=-32;
sine[19336]=-32;
sine[19337]=-32;
sine[19338]=-32;
sine[19339]=-32;
sine[19340]=-31;
sine[19341]=-31;
sine[19342]=-31;
sine[19343]=-31;
sine[19344]=-31;
sine[19345]=-31;
sine[19346]=-31;
sine[19347]=-31;
sine[19348]=-31;
sine[19349]=-31;
sine[19350]=-31;
sine[19351]=-31;
sine[19352]=-31;
sine[19353]=-31;
sine[19354]=-31;
sine[19355]=-31;
sine[19356]=-31;
sine[19357]=-31;
sine[19358]=-31;
sine[19359]=-31;
sine[19360]=-31;
sine[19361]=-31;
sine[19362]=-30;
sine[19363]=-30;
sine[19364]=-30;
sine[19365]=-30;
sine[19366]=-30;
sine[19367]=-30;
sine[19368]=-30;
sine[19369]=-30;
sine[19370]=-30;
sine[19371]=-30;
sine[19372]=-30;
sine[19373]=-30;
sine[19374]=-30;
sine[19375]=-30;
sine[19376]=-30;
sine[19377]=-30;
sine[19378]=-30;
sine[19379]=-30;
sine[19380]=-30;
sine[19381]=-30;
sine[19382]=-30;
sine[19383]=-30;
sine[19384]=-29;
sine[19385]=-29;
sine[19386]=-29;
sine[19387]=-29;
sine[19388]=-29;
sine[19389]=-29;
sine[19390]=-29;
sine[19391]=-29;
sine[19392]=-29;
sine[19393]=-29;
sine[19394]=-29;
sine[19395]=-29;
sine[19396]=-29;
sine[19397]=-29;
sine[19398]=-29;
sine[19399]=-29;
sine[19400]=-29;
sine[19401]=-29;
sine[19402]=-29;
sine[19403]=-29;
sine[19404]=-29;
sine[19405]=-29;
sine[19406]=-28;
sine[19407]=-28;
sine[19408]=-28;
sine[19409]=-28;
sine[19410]=-28;
sine[19411]=-28;
sine[19412]=-28;
sine[19413]=-28;
sine[19414]=-28;
sine[19415]=-28;
sine[19416]=-28;
sine[19417]=-28;
sine[19418]=-28;
sine[19419]=-28;
sine[19420]=-28;
sine[19421]=-28;
sine[19422]=-28;
sine[19423]=-28;
sine[19424]=-28;
sine[19425]=-28;
sine[19426]=-28;
sine[19427]=-28;
sine[19428]=-27;
sine[19429]=-27;
sine[19430]=-27;
sine[19431]=-27;
sine[19432]=-27;
sine[19433]=-27;
sine[19434]=-27;
sine[19435]=-27;
sine[19436]=-27;
sine[19437]=-27;
sine[19438]=-27;
sine[19439]=-27;
sine[19440]=-27;
sine[19441]=-27;
sine[19442]=-27;
sine[19443]=-27;
sine[19444]=-27;
sine[19445]=-27;
sine[19446]=-27;
sine[19447]=-27;
sine[19448]=-27;
sine[19449]=-27;
sine[19450]=-26;
sine[19451]=-26;
sine[19452]=-26;
sine[19453]=-26;
sine[19454]=-26;
sine[19455]=-26;
sine[19456]=-26;
sine[19457]=-26;
sine[19458]=-26;
sine[19459]=-26;
sine[19460]=-26;
sine[19461]=-26;
sine[19462]=-26;
sine[19463]=-26;
sine[19464]=-26;
sine[19465]=-26;
sine[19466]=-26;
sine[19467]=-26;
sine[19468]=-26;
sine[19469]=-26;
sine[19470]=-26;
sine[19471]=-25;
sine[19472]=-25;
sine[19473]=-25;
sine[19474]=-25;
sine[19475]=-25;
sine[19476]=-25;
sine[19477]=-25;
sine[19478]=-25;
sine[19479]=-25;
sine[19480]=-25;
sine[19481]=-25;
sine[19482]=-25;
sine[19483]=-25;
sine[19484]=-25;
sine[19485]=-25;
sine[19486]=-25;
sine[19487]=-25;
sine[19488]=-25;
sine[19489]=-25;
sine[19490]=-25;
sine[19491]=-25;
sine[19492]=-25;
sine[19493]=-24;
sine[19494]=-24;
sine[19495]=-24;
sine[19496]=-24;
sine[19497]=-24;
sine[19498]=-24;
sine[19499]=-24;
sine[19500]=-24;
sine[19501]=-24;
sine[19502]=-24;
sine[19503]=-24;
sine[19504]=-24;
sine[19505]=-24;
sine[19506]=-24;
sine[19507]=-24;
sine[19508]=-24;
sine[19509]=-24;
sine[19510]=-24;
sine[19511]=-24;
sine[19512]=-24;
sine[19513]=-24;
sine[19514]=-23;
sine[19515]=-23;
sine[19516]=-23;
sine[19517]=-23;
sine[19518]=-23;
sine[19519]=-23;
sine[19520]=-23;
sine[19521]=-23;
sine[19522]=-23;
sine[19523]=-23;
sine[19524]=-23;
sine[19525]=-23;
sine[19526]=-23;
sine[19527]=-23;
sine[19528]=-23;
sine[19529]=-23;
sine[19530]=-23;
sine[19531]=-23;
sine[19532]=-23;
sine[19533]=-23;
sine[19534]=-23;
sine[19535]=-23;
sine[19536]=-22;
sine[19537]=-22;
sine[19538]=-22;
sine[19539]=-22;
sine[19540]=-22;
sine[19541]=-22;
sine[19542]=-22;
sine[19543]=-22;
sine[19544]=-22;
sine[19545]=-22;
sine[19546]=-22;
sine[19547]=-22;
sine[19548]=-22;
sine[19549]=-22;
sine[19550]=-22;
sine[19551]=-22;
sine[19552]=-22;
sine[19553]=-22;
sine[19554]=-22;
sine[19555]=-22;
sine[19556]=-22;
sine[19557]=-21;
sine[19558]=-21;
sine[19559]=-21;
sine[19560]=-21;
sine[19561]=-21;
sine[19562]=-21;
sine[19563]=-21;
sine[19564]=-21;
sine[19565]=-21;
sine[19566]=-21;
sine[19567]=-21;
sine[19568]=-21;
sine[19569]=-21;
sine[19570]=-21;
sine[19571]=-21;
sine[19572]=-21;
sine[19573]=-21;
sine[19574]=-21;
sine[19575]=-21;
sine[19576]=-21;
sine[19577]=-21;
sine[19578]=-20;
sine[19579]=-20;
sine[19580]=-20;
sine[19581]=-20;
sine[19582]=-20;
sine[19583]=-20;
sine[19584]=-20;
sine[19585]=-20;
sine[19586]=-20;
sine[19587]=-20;
sine[19588]=-20;
sine[19589]=-20;
sine[19590]=-20;
sine[19591]=-20;
sine[19592]=-20;
sine[19593]=-20;
sine[19594]=-20;
sine[19595]=-20;
sine[19596]=-20;
sine[19597]=-20;
sine[19598]=-20;
sine[19599]=-19;
sine[19600]=-19;
sine[19601]=-19;
sine[19602]=-19;
sine[19603]=-19;
sine[19604]=-19;
sine[19605]=-19;
sine[19606]=-19;
sine[19607]=-19;
sine[19608]=-19;
sine[19609]=-19;
sine[19610]=-19;
sine[19611]=-19;
sine[19612]=-19;
sine[19613]=-19;
sine[19614]=-19;
sine[19615]=-19;
sine[19616]=-19;
sine[19617]=-19;
sine[19618]=-19;
sine[19619]=-19;
sine[19620]=-18;
sine[19621]=-18;
sine[19622]=-18;
sine[19623]=-18;
sine[19624]=-18;
sine[19625]=-18;
sine[19626]=-18;
sine[19627]=-18;
sine[19628]=-18;
sine[19629]=-18;
sine[19630]=-18;
sine[19631]=-18;
sine[19632]=-18;
sine[19633]=-18;
sine[19634]=-18;
sine[19635]=-18;
sine[19636]=-18;
sine[19637]=-18;
sine[19638]=-18;
sine[19639]=-18;
sine[19640]=-18;
sine[19641]=-17;
sine[19642]=-17;
sine[19643]=-17;
sine[19644]=-17;
sine[19645]=-17;
sine[19646]=-17;
sine[19647]=-17;
sine[19648]=-17;
sine[19649]=-17;
sine[19650]=-17;
sine[19651]=-17;
sine[19652]=-17;
sine[19653]=-17;
sine[19654]=-17;
sine[19655]=-17;
sine[19656]=-17;
sine[19657]=-17;
sine[19658]=-17;
sine[19659]=-17;
sine[19660]=-17;
sine[19661]=-17;
sine[19662]=-16;
sine[19663]=-16;
sine[19664]=-16;
sine[19665]=-16;
sine[19666]=-16;
sine[19667]=-16;
sine[19668]=-16;
sine[19669]=-16;
sine[19670]=-16;
sine[19671]=-16;
sine[19672]=-16;
sine[19673]=-16;
sine[19674]=-16;
sine[19675]=-16;
sine[19676]=-16;
sine[19677]=-16;
sine[19678]=-16;
sine[19679]=-16;
sine[19680]=-16;
sine[19681]=-16;
sine[19682]=-16;
sine[19683]=-15;
sine[19684]=-15;
sine[19685]=-15;
sine[19686]=-15;
sine[19687]=-15;
sine[19688]=-15;
sine[19689]=-15;
sine[19690]=-15;
sine[19691]=-15;
sine[19692]=-15;
sine[19693]=-15;
sine[19694]=-15;
sine[19695]=-15;
sine[19696]=-15;
sine[19697]=-15;
sine[19698]=-15;
sine[19699]=-15;
sine[19700]=-15;
sine[19701]=-15;
sine[19702]=-15;
sine[19703]=-14;
sine[19704]=-14;
sine[19705]=-14;
sine[19706]=-14;
sine[19707]=-14;
sine[19708]=-14;
sine[19709]=-14;
sine[19710]=-14;
sine[19711]=-14;
sine[19712]=-14;
sine[19713]=-14;
sine[19714]=-14;
sine[19715]=-14;
sine[19716]=-14;
sine[19717]=-14;
sine[19718]=-14;
sine[19719]=-14;
sine[19720]=-14;
sine[19721]=-14;
sine[19722]=-14;
sine[19723]=-14;
sine[19724]=-13;
sine[19725]=-13;
sine[19726]=-13;
sine[19727]=-13;
sine[19728]=-13;
sine[19729]=-13;
sine[19730]=-13;
sine[19731]=-13;
sine[19732]=-13;
sine[19733]=-13;
sine[19734]=-13;
sine[19735]=-13;
sine[19736]=-13;
sine[19737]=-13;
sine[19738]=-13;
sine[19739]=-13;
sine[19740]=-13;
sine[19741]=-13;
sine[19742]=-13;
sine[19743]=-13;
sine[19744]=-13;
sine[19745]=-12;
sine[19746]=-12;
sine[19747]=-12;
sine[19748]=-12;
sine[19749]=-12;
sine[19750]=-12;
sine[19751]=-12;
sine[19752]=-12;
sine[19753]=-12;
sine[19754]=-12;
sine[19755]=-12;
sine[19756]=-12;
sine[19757]=-12;
sine[19758]=-12;
sine[19759]=-12;
sine[19760]=-12;
sine[19761]=-12;
sine[19762]=-12;
sine[19763]=-12;
sine[19764]=-12;
sine[19765]=-11;
sine[19766]=-11;
sine[19767]=-11;
sine[19768]=-11;
sine[19769]=-11;
sine[19770]=-11;
sine[19771]=-11;
sine[19772]=-11;
sine[19773]=-11;
sine[19774]=-11;
sine[19775]=-11;
sine[19776]=-11;
sine[19777]=-11;
sine[19778]=-11;
sine[19779]=-11;
sine[19780]=-11;
sine[19781]=-11;
sine[19782]=-11;
sine[19783]=-11;
sine[19784]=-11;
sine[19785]=-11;
sine[19786]=-10;
sine[19787]=-10;
sine[19788]=-10;
sine[19789]=-10;
sine[19790]=-10;
sine[19791]=-10;
sine[19792]=-10;
sine[19793]=-10;
sine[19794]=-10;
sine[19795]=-10;
sine[19796]=-10;
sine[19797]=-10;
sine[19798]=-10;
sine[19799]=-10;
sine[19800]=-10;
sine[19801]=-10;
sine[19802]=-10;
sine[19803]=-10;
sine[19804]=-10;
sine[19805]=-10;
sine[19806]=-9;
sine[19807]=-9;
sine[19808]=-9;
sine[19809]=-9;
sine[19810]=-9;
sine[19811]=-9;
sine[19812]=-9;
sine[19813]=-9;
sine[19814]=-9;
sine[19815]=-9;
sine[19816]=-9;
sine[19817]=-9;
sine[19818]=-9;
sine[19819]=-9;
sine[19820]=-9;
sine[19821]=-9;
sine[19822]=-9;
sine[19823]=-9;
sine[19824]=-9;
sine[19825]=-9;
sine[19826]=-9;
sine[19827]=-8;
sine[19828]=-8;
sine[19829]=-8;
sine[19830]=-8;
sine[19831]=-8;
sine[19832]=-8;
sine[19833]=-8;
sine[19834]=-8;
sine[19835]=-8;
sine[19836]=-8;
sine[19837]=-8;
sine[19838]=-8;
sine[19839]=-8;
sine[19840]=-8;
sine[19841]=-8;
sine[19842]=-8;
sine[19843]=-8;
sine[19844]=-8;
sine[19845]=-8;
sine[19846]=-8;
sine[19847]=-7;
sine[19848]=-7;
sine[19849]=-7;
sine[19850]=-7;
sine[19851]=-7;
sine[19852]=-7;
sine[19853]=-7;
sine[19854]=-7;
sine[19855]=-7;
sine[19856]=-7;
sine[19857]=-7;
sine[19858]=-7;
sine[19859]=-7;
sine[19860]=-7;
sine[19861]=-7;
sine[19862]=-7;
sine[19863]=-7;
sine[19864]=-7;
sine[19865]=-7;
sine[19866]=-7;
sine[19867]=-7;
sine[19868]=-6;
sine[19869]=-6;
sine[19870]=-6;
sine[19871]=-6;
sine[19872]=-6;
sine[19873]=-6;
sine[19874]=-6;
sine[19875]=-6;
sine[19876]=-6;
sine[19877]=-6;
sine[19878]=-6;
sine[19879]=-6;
sine[19880]=-6;
sine[19881]=-6;
sine[19882]=-6;
sine[19883]=-6;
sine[19884]=-6;
sine[19885]=-6;
sine[19886]=-6;
sine[19887]=-6;
sine[19888]=-5;
sine[19889]=-5;
sine[19890]=-5;
sine[19891]=-5;
sine[19892]=-5;
sine[19893]=-5;
sine[19894]=-5;
sine[19895]=-5;
sine[19896]=-5;
sine[19897]=-5;
sine[19898]=-5;
sine[19899]=-5;
sine[19900]=-5;
sine[19901]=-5;
sine[19902]=-5;
sine[19903]=-5;
sine[19904]=-5;
sine[19905]=-5;
sine[19906]=-5;
sine[19907]=-5;
sine[19908]=-5;
sine[19909]=-4;
sine[19910]=-4;
sine[19911]=-4;
sine[19912]=-4;
sine[19913]=-4;
sine[19914]=-4;
sine[19915]=-4;
sine[19916]=-4;
sine[19917]=-4;
sine[19918]=-4;
sine[19919]=-4;
sine[19920]=-4;
sine[19921]=-4;
sine[19922]=-4;
sine[19923]=-4;
sine[19924]=-4;
sine[19925]=-4;
sine[19926]=-4;
sine[19927]=-4;
sine[19928]=-4;
sine[19929]=-3;
sine[19930]=-3;
sine[19931]=-3;
sine[19932]=-3;
sine[19933]=-3;
sine[19934]=-3;
sine[19935]=-3;
sine[19936]=-3;
sine[19937]=-3;
sine[19938]=-3;
sine[19939]=-3;
sine[19940]=-3;
sine[19941]=-3;
sine[19942]=-3;
sine[19943]=-3;
sine[19944]=-3;
sine[19945]=-3;
sine[19946]=-3;
sine[19947]=-3;
sine[19948]=-3;
sine[19949]=-3;
sine[19950]=-2;
sine[19951]=-2;
sine[19952]=-2;
sine[19953]=-2;
sine[19954]=-2;
sine[19955]=-2;
sine[19956]=-2;
sine[19957]=-2;
sine[19958]=-2;
sine[19959]=-2;
sine[19960]=-2;
sine[19961]=-2;
sine[19962]=-2;
sine[19963]=-2;
sine[19964]=-2;
sine[19965]=-2;
sine[19966]=-2;
sine[19967]=-2;
sine[19968]=-2;
sine[19969]=-2;
sine[19970]=-1;
sine[19971]=-1;
sine[19972]=-1;
sine[19973]=-1;
sine[19974]=-1;
sine[19975]=-1;
sine[19976]=-1;
sine[19977]=-1;
sine[19978]=-1;
sine[19979]=-1;
sine[19980]=-1;
sine[19981]=-1;
sine[19982]=-1;
sine[19983]=-1;
sine[19984]=-1;
sine[19985]=-1;
sine[19986]=-1;
sine[19987]=-1;
sine[19988]=-1;
sine[19989]=-1;
sine[19990]=0;
sine[19991]=0;
sine[19992]=0;
sine[19993]=0;
sine[19994]=0;
sine[19995]=0;
sine[19996]=0;
sine[19997]=0;
sine[19998]=0;
sine[19999]=0;
sine[20000]=0;
sine[20001]=0;
sine[20002]=0;
sine[20003]=0;
sine[20004]=0;
sine[20005]=0;
sine[20006]=0;
sine[20007]=0;
sine[20008]=0;
sine[20009]=0;
sine[20010]=0;
sine[20011]=1;
sine[20012]=1;
sine[20013]=1;
sine[20014]=1;
sine[20015]=1;
sine[20016]=1;
sine[20017]=1;
sine[20018]=1;
sine[20019]=1;
sine[20020]=1;
sine[20021]=1;
sine[20022]=1;
sine[20023]=1;
sine[20024]=1;
sine[20025]=1;
sine[20026]=1;
sine[20027]=1;
sine[20028]=1;
sine[20029]=1;
sine[20030]=1;
sine[20031]=2;
sine[20032]=2;
sine[20033]=2;
sine[20034]=2;
sine[20035]=2;
sine[20036]=2;
sine[20037]=2;
sine[20038]=2;
sine[20039]=2;
sine[20040]=2;
sine[20041]=2;
sine[20042]=2;
sine[20043]=2;
sine[20044]=2;
sine[20045]=2;
sine[20046]=2;
sine[20047]=2;
sine[20048]=2;
sine[20049]=2;
sine[20050]=2;
sine[20051]=3;
sine[20052]=3;
sine[20053]=3;
sine[20054]=3;
sine[20055]=3;
sine[20056]=3;
sine[20057]=3;
sine[20058]=3;
sine[20059]=3;
sine[20060]=3;
sine[20061]=3;
sine[20062]=3;
sine[20063]=3;
sine[20064]=3;
sine[20065]=3;
sine[20066]=3;
sine[20067]=3;
sine[20068]=3;
sine[20069]=3;
sine[20070]=3;
sine[20071]=3;
sine[20072]=4;
sine[20073]=4;
sine[20074]=4;
sine[20075]=4;
sine[20076]=4;
sine[20077]=4;
sine[20078]=4;
sine[20079]=4;
sine[20080]=4;
sine[20081]=4;
sine[20082]=4;
sine[20083]=4;
sine[20084]=4;
sine[20085]=4;
sine[20086]=4;
sine[20087]=4;
sine[20088]=4;
sine[20089]=4;
sine[20090]=4;
sine[20091]=4;
sine[20092]=5;
sine[20093]=5;
sine[20094]=5;
sine[20095]=5;
sine[20096]=5;
sine[20097]=5;
sine[20098]=5;
sine[20099]=5;
sine[20100]=5;
sine[20101]=5;
sine[20102]=5;
sine[20103]=5;
sine[20104]=5;
sine[20105]=5;
sine[20106]=5;
sine[20107]=5;
sine[20108]=5;
sine[20109]=5;
sine[20110]=5;
sine[20111]=5;
sine[20112]=5;
sine[20113]=6;
sine[20114]=6;
sine[20115]=6;
sine[20116]=6;
sine[20117]=6;
sine[20118]=6;
sine[20119]=6;
sine[20120]=6;
sine[20121]=6;
sine[20122]=6;
sine[20123]=6;
sine[20124]=6;
sine[20125]=6;
sine[20126]=6;
sine[20127]=6;
sine[20128]=6;
sine[20129]=6;
sine[20130]=6;
sine[20131]=6;
sine[20132]=6;
sine[20133]=7;
sine[20134]=7;
sine[20135]=7;
sine[20136]=7;
sine[20137]=7;
sine[20138]=7;
sine[20139]=7;
sine[20140]=7;
sine[20141]=7;
sine[20142]=7;
sine[20143]=7;
sine[20144]=7;
sine[20145]=7;
sine[20146]=7;
sine[20147]=7;
sine[20148]=7;
sine[20149]=7;
sine[20150]=7;
sine[20151]=7;
sine[20152]=7;
sine[20153]=7;
sine[20154]=8;
sine[20155]=8;
sine[20156]=8;
sine[20157]=8;
sine[20158]=8;
sine[20159]=8;
sine[20160]=8;
sine[20161]=8;
sine[20162]=8;
sine[20163]=8;
sine[20164]=8;
sine[20165]=8;
sine[20166]=8;
sine[20167]=8;
sine[20168]=8;
sine[20169]=8;
sine[20170]=8;
sine[20171]=8;
sine[20172]=8;
sine[20173]=8;
sine[20174]=9;
sine[20175]=9;
sine[20176]=9;
sine[20177]=9;
sine[20178]=9;
sine[20179]=9;
sine[20180]=9;
sine[20181]=9;
sine[20182]=9;
sine[20183]=9;
sine[20184]=9;
sine[20185]=9;
sine[20186]=9;
sine[20187]=9;
sine[20188]=9;
sine[20189]=9;
sine[20190]=9;
sine[20191]=9;
sine[20192]=9;
sine[20193]=9;
sine[20194]=9;
sine[20195]=10;
sine[20196]=10;
sine[20197]=10;
sine[20198]=10;
sine[20199]=10;
sine[20200]=10;
sine[20201]=10;
sine[20202]=10;
sine[20203]=10;
sine[20204]=10;
sine[20205]=10;
sine[20206]=10;
sine[20207]=10;
sine[20208]=10;
sine[20209]=10;
sine[20210]=10;
sine[20211]=10;
sine[20212]=10;
sine[20213]=10;
sine[20214]=10;
sine[20215]=11;
sine[20216]=11;
sine[20217]=11;
sine[20218]=11;
sine[20219]=11;
sine[20220]=11;
sine[20221]=11;
sine[20222]=11;
sine[20223]=11;
sine[20224]=11;
sine[20225]=11;
sine[20226]=11;
sine[20227]=11;
sine[20228]=11;
sine[20229]=11;
sine[20230]=11;
sine[20231]=11;
sine[20232]=11;
sine[20233]=11;
sine[20234]=11;
sine[20235]=11;
sine[20236]=12;
sine[20237]=12;
sine[20238]=12;
sine[20239]=12;
sine[20240]=12;
sine[20241]=12;
sine[20242]=12;
sine[20243]=12;
sine[20244]=12;
sine[20245]=12;
sine[20246]=12;
sine[20247]=12;
sine[20248]=12;
sine[20249]=12;
sine[20250]=12;
sine[20251]=12;
sine[20252]=12;
sine[20253]=12;
sine[20254]=12;
sine[20255]=12;
sine[20256]=13;
sine[20257]=13;
sine[20258]=13;
sine[20259]=13;
sine[20260]=13;
sine[20261]=13;
sine[20262]=13;
sine[20263]=13;
sine[20264]=13;
sine[20265]=13;
sine[20266]=13;
sine[20267]=13;
sine[20268]=13;
sine[20269]=13;
sine[20270]=13;
sine[20271]=13;
sine[20272]=13;
sine[20273]=13;
sine[20274]=13;
sine[20275]=13;
sine[20276]=13;
sine[20277]=14;
sine[20278]=14;
sine[20279]=14;
sine[20280]=14;
sine[20281]=14;
sine[20282]=14;
sine[20283]=14;
sine[20284]=14;
sine[20285]=14;
sine[20286]=14;
sine[20287]=14;
sine[20288]=14;
sine[20289]=14;
sine[20290]=14;
sine[20291]=14;
sine[20292]=14;
sine[20293]=14;
sine[20294]=14;
sine[20295]=14;
sine[20296]=14;
sine[20297]=14;
sine[20298]=15;
sine[20299]=15;
sine[20300]=15;
sine[20301]=15;
sine[20302]=15;
sine[20303]=15;
sine[20304]=15;
sine[20305]=15;
sine[20306]=15;
sine[20307]=15;
sine[20308]=15;
sine[20309]=15;
sine[20310]=15;
sine[20311]=15;
sine[20312]=15;
sine[20313]=15;
sine[20314]=15;
sine[20315]=15;
sine[20316]=15;
sine[20317]=15;
sine[20318]=16;
sine[20319]=16;
sine[20320]=16;
sine[20321]=16;
sine[20322]=16;
sine[20323]=16;
sine[20324]=16;
sine[20325]=16;
sine[20326]=16;
sine[20327]=16;
sine[20328]=16;
sine[20329]=16;
sine[20330]=16;
sine[20331]=16;
sine[20332]=16;
sine[20333]=16;
sine[20334]=16;
sine[20335]=16;
sine[20336]=16;
sine[20337]=16;
sine[20338]=16;
sine[20339]=17;
sine[20340]=17;
sine[20341]=17;
sine[20342]=17;
sine[20343]=17;
sine[20344]=17;
sine[20345]=17;
sine[20346]=17;
sine[20347]=17;
sine[20348]=17;
sine[20349]=17;
sine[20350]=17;
sine[20351]=17;
sine[20352]=17;
sine[20353]=17;
sine[20354]=17;
sine[20355]=17;
sine[20356]=17;
sine[20357]=17;
sine[20358]=17;
sine[20359]=17;
sine[20360]=18;
sine[20361]=18;
sine[20362]=18;
sine[20363]=18;
sine[20364]=18;
sine[20365]=18;
sine[20366]=18;
sine[20367]=18;
sine[20368]=18;
sine[20369]=18;
sine[20370]=18;
sine[20371]=18;
sine[20372]=18;
sine[20373]=18;
sine[20374]=18;
sine[20375]=18;
sine[20376]=18;
sine[20377]=18;
sine[20378]=18;
sine[20379]=18;
sine[20380]=18;
sine[20381]=19;
sine[20382]=19;
sine[20383]=19;
sine[20384]=19;
sine[20385]=19;
sine[20386]=19;
sine[20387]=19;
sine[20388]=19;
sine[20389]=19;
sine[20390]=19;
sine[20391]=19;
sine[20392]=19;
sine[20393]=19;
sine[20394]=19;
sine[20395]=19;
sine[20396]=19;
sine[20397]=19;
sine[20398]=19;
sine[20399]=19;
sine[20400]=19;
sine[20401]=19;
sine[20402]=20;
sine[20403]=20;
sine[20404]=20;
sine[20405]=20;
sine[20406]=20;
sine[20407]=20;
sine[20408]=20;
sine[20409]=20;
sine[20410]=20;
sine[20411]=20;
sine[20412]=20;
sine[20413]=20;
sine[20414]=20;
sine[20415]=20;
sine[20416]=20;
sine[20417]=20;
sine[20418]=20;
sine[20419]=20;
sine[20420]=20;
sine[20421]=20;
sine[20422]=20;
sine[20423]=21;
sine[20424]=21;
sine[20425]=21;
sine[20426]=21;
sine[20427]=21;
sine[20428]=21;
sine[20429]=21;
sine[20430]=21;
sine[20431]=21;
sine[20432]=21;
sine[20433]=21;
sine[20434]=21;
sine[20435]=21;
sine[20436]=21;
sine[20437]=21;
sine[20438]=21;
sine[20439]=21;
sine[20440]=21;
sine[20441]=21;
sine[20442]=21;
sine[20443]=21;
sine[20444]=22;
sine[20445]=22;
sine[20446]=22;
sine[20447]=22;
sine[20448]=22;
sine[20449]=22;
sine[20450]=22;
sine[20451]=22;
sine[20452]=22;
sine[20453]=22;
sine[20454]=22;
sine[20455]=22;
sine[20456]=22;
sine[20457]=22;
sine[20458]=22;
sine[20459]=22;
sine[20460]=22;
sine[20461]=22;
sine[20462]=22;
sine[20463]=22;
sine[20464]=22;
sine[20465]=23;
sine[20466]=23;
sine[20467]=23;
sine[20468]=23;
sine[20469]=23;
sine[20470]=23;
sine[20471]=23;
sine[20472]=23;
sine[20473]=23;
sine[20474]=23;
sine[20475]=23;
sine[20476]=23;
sine[20477]=23;
sine[20478]=23;
sine[20479]=23;
sine[20480]=23;
sine[20481]=23;
sine[20482]=23;
sine[20483]=23;
sine[20484]=23;
sine[20485]=23;
sine[20486]=23;
sine[20487]=24;
sine[20488]=24;
sine[20489]=24;
sine[20490]=24;
sine[20491]=24;
sine[20492]=24;
sine[20493]=24;
sine[20494]=24;
sine[20495]=24;
sine[20496]=24;
sine[20497]=24;
sine[20498]=24;
sine[20499]=24;
sine[20500]=24;
sine[20501]=24;
sine[20502]=24;
sine[20503]=24;
sine[20504]=24;
sine[20505]=24;
sine[20506]=24;
sine[20507]=24;
sine[20508]=25;
sine[20509]=25;
sine[20510]=25;
sine[20511]=25;
sine[20512]=25;
sine[20513]=25;
sine[20514]=25;
sine[20515]=25;
sine[20516]=25;
sine[20517]=25;
sine[20518]=25;
sine[20519]=25;
sine[20520]=25;
sine[20521]=25;
sine[20522]=25;
sine[20523]=25;
sine[20524]=25;
sine[20525]=25;
sine[20526]=25;
sine[20527]=25;
sine[20528]=25;
sine[20529]=25;
sine[20530]=26;
sine[20531]=26;
sine[20532]=26;
sine[20533]=26;
sine[20534]=26;
sine[20535]=26;
sine[20536]=26;
sine[20537]=26;
sine[20538]=26;
sine[20539]=26;
sine[20540]=26;
sine[20541]=26;
sine[20542]=26;
sine[20543]=26;
sine[20544]=26;
sine[20545]=26;
sine[20546]=26;
sine[20547]=26;
sine[20548]=26;
sine[20549]=26;
sine[20550]=26;
sine[20551]=27;
sine[20552]=27;
sine[20553]=27;
sine[20554]=27;
sine[20555]=27;
sine[20556]=27;
sine[20557]=27;
sine[20558]=27;
sine[20559]=27;
sine[20560]=27;
sine[20561]=27;
sine[20562]=27;
sine[20563]=27;
sine[20564]=27;
sine[20565]=27;
sine[20566]=27;
sine[20567]=27;
sine[20568]=27;
sine[20569]=27;
sine[20570]=27;
sine[20571]=27;
sine[20572]=27;
sine[20573]=28;
sine[20574]=28;
sine[20575]=28;
sine[20576]=28;
sine[20577]=28;
sine[20578]=28;
sine[20579]=28;
sine[20580]=28;
sine[20581]=28;
sine[20582]=28;
sine[20583]=28;
sine[20584]=28;
sine[20585]=28;
sine[20586]=28;
sine[20587]=28;
sine[20588]=28;
sine[20589]=28;
sine[20590]=28;
sine[20591]=28;
sine[20592]=28;
sine[20593]=28;
sine[20594]=28;
sine[20595]=29;
sine[20596]=29;
sine[20597]=29;
sine[20598]=29;
sine[20599]=29;
sine[20600]=29;
sine[20601]=29;
sine[20602]=29;
sine[20603]=29;
sine[20604]=29;
sine[20605]=29;
sine[20606]=29;
sine[20607]=29;
sine[20608]=29;
sine[20609]=29;
sine[20610]=29;
sine[20611]=29;
sine[20612]=29;
sine[20613]=29;
sine[20614]=29;
sine[20615]=29;
sine[20616]=29;
sine[20617]=30;
sine[20618]=30;
sine[20619]=30;
sine[20620]=30;
sine[20621]=30;
sine[20622]=30;
sine[20623]=30;
sine[20624]=30;
sine[20625]=30;
sine[20626]=30;
sine[20627]=30;
sine[20628]=30;
sine[20629]=30;
sine[20630]=30;
sine[20631]=30;
sine[20632]=30;
sine[20633]=30;
sine[20634]=30;
sine[20635]=30;
sine[20636]=30;
sine[20637]=30;
sine[20638]=30;
sine[20639]=31;
sine[20640]=31;
sine[20641]=31;
sine[20642]=31;
sine[20643]=31;
sine[20644]=31;
sine[20645]=31;
sine[20646]=31;
sine[20647]=31;
sine[20648]=31;
sine[20649]=31;
sine[20650]=31;
sine[20651]=31;
sine[20652]=31;
sine[20653]=31;
sine[20654]=31;
sine[20655]=31;
sine[20656]=31;
sine[20657]=31;
sine[20658]=31;
sine[20659]=31;
sine[20660]=31;
sine[20661]=32;
sine[20662]=32;
sine[20663]=32;
sine[20664]=32;
sine[20665]=32;
sine[20666]=32;
sine[20667]=32;
sine[20668]=32;
sine[20669]=32;
sine[20670]=32;
sine[20671]=32;
sine[20672]=32;
sine[20673]=32;
sine[20674]=32;
sine[20675]=32;
sine[20676]=32;
sine[20677]=32;
sine[20678]=32;
sine[20679]=32;
sine[20680]=32;
sine[20681]=32;
sine[20682]=32;
sine[20683]=33;
sine[20684]=33;
sine[20685]=33;
sine[20686]=33;
sine[20687]=33;
sine[20688]=33;
sine[20689]=33;
sine[20690]=33;
sine[20691]=33;
sine[20692]=33;
sine[20693]=33;
sine[20694]=33;
sine[20695]=33;
sine[20696]=33;
sine[20697]=33;
sine[20698]=33;
sine[20699]=33;
sine[20700]=33;
sine[20701]=33;
sine[20702]=33;
sine[20703]=33;
sine[20704]=33;
sine[20705]=33;
sine[20706]=34;
sine[20707]=34;
sine[20708]=34;
sine[20709]=34;
sine[20710]=34;
sine[20711]=34;
sine[20712]=34;
sine[20713]=34;
sine[20714]=34;
sine[20715]=34;
sine[20716]=34;
sine[20717]=34;
sine[20718]=34;
sine[20719]=34;
sine[20720]=34;
sine[20721]=34;
sine[20722]=34;
sine[20723]=34;
sine[20724]=34;
sine[20725]=34;
sine[20726]=34;
sine[20727]=34;
sine[20728]=35;
sine[20729]=35;
sine[20730]=35;
sine[20731]=35;
sine[20732]=35;
sine[20733]=35;
sine[20734]=35;
sine[20735]=35;
sine[20736]=35;
sine[20737]=35;
sine[20738]=35;
sine[20739]=35;
sine[20740]=35;
sine[20741]=35;
sine[20742]=35;
sine[20743]=35;
sine[20744]=35;
sine[20745]=35;
sine[20746]=35;
sine[20747]=35;
sine[20748]=35;
sine[20749]=35;
sine[20750]=35;
sine[20751]=36;
sine[20752]=36;
sine[20753]=36;
sine[20754]=36;
sine[20755]=36;
sine[20756]=36;
sine[20757]=36;
sine[20758]=36;
sine[20759]=36;
sine[20760]=36;
sine[20761]=36;
sine[20762]=36;
sine[20763]=36;
sine[20764]=36;
sine[20765]=36;
sine[20766]=36;
sine[20767]=36;
sine[20768]=36;
sine[20769]=36;
sine[20770]=36;
sine[20771]=36;
sine[20772]=36;
sine[20773]=36;
sine[20774]=37;
sine[20775]=37;
sine[20776]=37;
sine[20777]=37;
sine[20778]=37;
sine[20779]=37;
sine[20780]=37;
sine[20781]=37;
sine[20782]=37;
sine[20783]=37;
sine[20784]=37;
sine[20785]=37;
sine[20786]=37;
sine[20787]=37;
sine[20788]=37;
sine[20789]=37;
sine[20790]=37;
sine[20791]=37;
sine[20792]=37;
sine[20793]=37;
sine[20794]=37;
sine[20795]=37;
sine[20796]=37;
sine[20797]=38;
sine[20798]=38;
sine[20799]=38;
sine[20800]=38;
sine[20801]=38;
sine[20802]=38;
sine[20803]=38;
sine[20804]=38;
sine[20805]=38;
sine[20806]=38;
sine[20807]=38;
sine[20808]=38;
sine[20809]=38;
sine[20810]=38;
sine[20811]=38;
sine[20812]=38;
sine[20813]=38;
sine[20814]=38;
sine[20815]=38;
sine[20816]=38;
sine[20817]=38;
sine[20818]=38;
sine[20819]=38;
sine[20820]=38;
sine[20821]=39;
sine[20822]=39;
sine[20823]=39;
sine[20824]=39;
sine[20825]=39;
sine[20826]=39;
sine[20827]=39;
sine[20828]=39;
sine[20829]=39;
sine[20830]=39;
sine[20831]=39;
sine[20832]=39;
sine[20833]=39;
sine[20834]=39;
sine[20835]=39;
sine[20836]=39;
sine[20837]=39;
sine[20838]=39;
sine[20839]=39;
sine[20840]=39;
sine[20841]=39;
sine[20842]=39;
sine[20843]=39;
sine[20844]=40;
sine[20845]=40;
sine[20846]=40;
sine[20847]=40;
sine[20848]=40;
sine[20849]=40;
sine[20850]=40;
sine[20851]=40;
sine[20852]=40;
sine[20853]=40;
sine[20854]=40;
sine[20855]=40;
sine[20856]=40;
sine[20857]=40;
sine[20858]=40;
sine[20859]=40;
sine[20860]=40;
sine[20861]=40;
sine[20862]=40;
sine[20863]=40;
sine[20864]=40;
sine[20865]=40;
sine[20866]=40;
sine[20867]=40;
sine[20868]=41;
sine[20869]=41;
sine[20870]=41;
sine[20871]=41;
sine[20872]=41;
sine[20873]=41;
sine[20874]=41;
sine[20875]=41;
sine[20876]=41;
sine[20877]=41;
sine[20878]=41;
sine[20879]=41;
sine[20880]=41;
sine[20881]=41;
sine[20882]=41;
sine[20883]=41;
sine[20884]=41;
sine[20885]=41;
sine[20886]=41;
sine[20887]=41;
sine[20888]=41;
sine[20889]=41;
sine[20890]=41;
sine[20891]=41;
sine[20892]=42;
sine[20893]=42;
sine[20894]=42;
sine[20895]=42;
sine[20896]=42;
sine[20897]=42;
sine[20898]=42;
sine[20899]=42;
sine[20900]=42;
sine[20901]=42;
sine[20902]=42;
sine[20903]=42;
sine[20904]=42;
sine[20905]=42;
sine[20906]=42;
sine[20907]=42;
sine[20908]=42;
sine[20909]=42;
sine[20910]=42;
sine[20911]=42;
sine[20912]=42;
sine[20913]=42;
sine[20914]=42;
sine[20915]=42;
sine[20916]=43;
sine[20917]=43;
sine[20918]=43;
sine[20919]=43;
sine[20920]=43;
sine[20921]=43;
sine[20922]=43;
sine[20923]=43;
sine[20924]=43;
sine[20925]=43;
sine[20926]=43;
sine[20927]=43;
sine[20928]=43;
sine[20929]=43;
sine[20930]=43;
sine[20931]=43;
sine[20932]=43;
sine[20933]=43;
sine[20934]=43;
sine[20935]=43;
sine[20936]=43;
sine[20937]=43;
sine[20938]=43;
sine[20939]=43;
sine[20940]=44;
sine[20941]=44;
sine[20942]=44;
sine[20943]=44;
sine[20944]=44;
sine[20945]=44;
sine[20946]=44;
sine[20947]=44;
sine[20948]=44;
sine[20949]=44;
sine[20950]=44;
sine[20951]=44;
sine[20952]=44;
sine[20953]=44;
sine[20954]=44;
sine[20955]=44;
sine[20956]=44;
sine[20957]=44;
sine[20958]=44;
sine[20959]=44;
sine[20960]=44;
sine[20961]=44;
sine[20962]=44;
sine[20963]=44;
sine[20964]=44;
sine[20965]=45;
sine[20966]=45;
sine[20967]=45;
sine[20968]=45;
sine[20969]=45;
sine[20970]=45;
sine[20971]=45;
sine[20972]=45;
sine[20973]=45;
sine[20974]=45;
sine[20975]=45;
sine[20976]=45;
sine[20977]=45;
sine[20978]=45;
sine[20979]=45;
sine[20980]=45;
sine[20981]=45;
sine[20982]=45;
sine[20983]=45;
sine[20984]=45;
sine[20985]=45;
sine[20986]=45;
sine[20987]=45;
sine[20988]=45;
sine[20989]=45;
sine[20990]=46;
sine[20991]=46;
sine[20992]=46;
sine[20993]=46;
sine[20994]=46;
sine[20995]=46;
sine[20996]=46;
sine[20997]=46;
sine[20998]=46;
sine[20999]=46;
sine[21000]=46;
sine[21001]=46;
sine[21002]=46;
sine[21003]=46;
sine[21004]=46;
sine[21005]=46;
sine[21006]=46;
sine[21007]=46;
sine[21008]=46;
sine[21009]=46;
sine[21010]=46;
sine[21011]=46;
sine[21012]=46;
sine[21013]=46;
sine[21014]=46;
sine[21015]=47;
sine[21016]=47;
sine[21017]=47;
sine[21018]=47;
sine[21019]=47;
sine[21020]=47;
sine[21021]=47;
sine[21022]=47;
sine[21023]=47;
sine[21024]=47;
sine[21025]=47;
sine[21026]=47;
sine[21027]=47;
sine[21028]=47;
sine[21029]=47;
sine[21030]=47;
sine[21031]=47;
sine[21032]=47;
sine[21033]=47;
sine[21034]=47;
sine[21035]=47;
sine[21036]=47;
sine[21037]=47;
sine[21038]=47;
sine[21039]=47;
sine[21040]=47;
sine[21041]=48;
sine[21042]=48;
sine[21043]=48;
sine[21044]=48;
sine[21045]=48;
sine[21046]=48;
sine[21047]=48;
sine[21048]=48;
sine[21049]=48;
sine[21050]=48;
sine[21051]=48;
sine[21052]=48;
sine[21053]=48;
sine[21054]=48;
sine[21055]=48;
sine[21056]=48;
sine[21057]=48;
sine[21058]=48;
sine[21059]=48;
sine[21060]=48;
sine[21061]=48;
sine[21062]=48;
sine[21063]=48;
sine[21064]=48;
sine[21065]=48;
sine[21066]=49;
sine[21067]=49;
sine[21068]=49;
sine[21069]=49;
sine[21070]=49;
sine[21071]=49;
sine[21072]=49;
sine[21073]=49;
sine[21074]=49;
sine[21075]=49;
sine[21076]=49;
sine[21077]=49;
sine[21078]=49;
sine[21079]=49;
sine[21080]=49;
sine[21081]=49;
sine[21082]=49;
sine[21083]=49;
sine[21084]=49;
sine[21085]=49;
sine[21086]=49;
sine[21087]=49;
sine[21088]=49;
sine[21089]=49;
sine[21090]=49;
sine[21091]=49;
sine[21092]=49;
sine[21093]=50;
sine[21094]=50;
sine[21095]=50;
sine[21096]=50;
sine[21097]=50;
sine[21098]=50;
sine[21099]=50;
sine[21100]=50;
sine[21101]=50;
sine[21102]=50;
sine[21103]=50;
sine[21104]=50;
sine[21105]=50;
sine[21106]=50;
sine[21107]=50;
sine[21108]=50;
sine[21109]=50;
sine[21110]=50;
sine[21111]=50;
sine[21112]=50;
sine[21113]=50;
sine[21114]=50;
sine[21115]=50;
sine[21116]=50;
sine[21117]=50;
sine[21118]=50;
sine[21119]=51;
sine[21120]=51;
sine[21121]=51;
sine[21122]=51;
sine[21123]=51;
sine[21124]=51;
sine[21125]=51;
sine[21126]=51;
sine[21127]=51;
sine[21128]=51;
sine[21129]=51;
sine[21130]=51;
sine[21131]=51;
sine[21132]=51;
sine[21133]=51;
sine[21134]=51;
sine[21135]=51;
sine[21136]=51;
sine[21137]=51;
sine[21138]=51;
sine[21139]=51;
sine[21140]=51;
sine[21141]=51;
sine[21142]=51;
sine[21143]=51;
sine[21144]=51;
sine[21145]=51;
sine[21146]=52;
sine[21147]=52;
sine[21148]=52;
sine[21149]=52;
sine[21150]=52;
sine[21151]=52;
sine[21152]=52;
sine[21153]=52;
sine[21154]=52;
sine[21155]=52;
sine[21156]=52;
sine[21157]=52;
sine[21158]=52;
sine[21159]=52;
sine[21160]=52;
sine[21161]=52;
sine[21162]=52;
sine[21163]=52;
sine[21164]=52;
sine[21165]=52;
sine[21166]=52;
sine[21167]=52;
sine[21168]=52;
sine[21169]=52;
sine[21170]=52;
sine[21171]=52;
sine[21172]=52;
sine[21173]=53;
sine[21174]=53;
sine[21175]=53;
sine[21176]=53;
sine[21177]=53;
sine[21178]=53;
sine[21179]=53;
sine[21180]=53;
sine[21181]=53;
sine[21182]=53;
sine[21183]=53;
sine[21184]=53;
sine[21185]=53;
sine[21186]=53;
sine[21187]=53;
sine[21188]=53;
sine[21189]=53;
sine[21190]=53;
sine[21191]=53;
sine[21192]=53;
sine[21193]=53;
sine[21194]=53;
sine[21195]=53;
sine[21196]=53;
sine[21197]=53;
sine[21198]=53;
sine[21199]=53;
sine[21200]=53;
sine[21201]=54;
sine[21202]=54;
sine[21203]=54;
sine[21204]=54;
sine[21205]=54;
sine[21206]=54;
sine[21207]=54;
sine[21208]=54;
sine[21209]=54;
sine[21210]=54;
sine[21211]=54;
sine[21212]=54;
sine[21213]=54;
sine[21214]=54;
sine[21215]=54;
sine[21216]=54;
sine[21217]=54;
sine[21218]=54;
sine[21219]=54;
sine[21220]=54;
sine[21221]=54;
sine[21222]=54;
sine[21223]=54;
sine[21224]=54;
sine[21225]=54;
sine[21226]=54;
sine[21227]=54;
sine[21228]=54;
sine[21229]=55;
sine[21230]=55;
sine[21231]=55;
sine[21232]=55;
sine[21233]=55;
sine[21234]=55;
sine[21235]=55;
sine[21236]=55;
sine[21237]=55;
sine[21238]=55;
sine[21239]=55;
sine[21240]=55;
sine[21241]=55;
sine[21242]=55;
sine[21243]=55;
sine[21244]=55;
sine[21245]=55;
sine[21246]=55;
sine[21247]=55;
sine[21248]=55;
sine[21249]=55;
sine[21250]=55;
sine[21251]=55;
sine[21252]=55;
sine[21253]=55;
sine[21254]=55;
sine[21255]=55;
sine[21256]=55;
sine[21257]=55;
sine[21258]=56;
sine[21259]=56;
sine[21260]=56;
sine[21261]=56;
sine[21262]=56;
sine[21263]=56;
sine[21264]=56;
sine[21265]=56;
sine[21266]=56;
sine[21267]=56;
sine[21268]=56;
sine[21269]=56;
sine[21270]=56;
sine[21271]=56;
sine[21272]=56;
sine[21273]=56;
sine[21274]=56;
sine[21275]=56;
sine[21276]=56;
sine[21277]=56;
sine[21278]=56;
sine[21279]=56;
sine[21280]=56;
sine[21281]=56;
sine[21282]=56;
sine[21283]=56;
sine[21284]=56;
sine[21285]=56;
sine[21286]=56;
sine[21287]=57;
sine[21288]=57;
sine[21289]=57;
sine[21290]=57;
sine[21291]=57;
sine[21292]=57;
sine[21293]=57;
sine[21294]=57;
sine[21295]=57;
sine[21296]=57;
sine[21297]=57;
sine[21298]=57;
sine[21299]=57;
sine[21300]=57;
sine[21301]=57;
sine[21302]=57;
sine[21303]=57;
sine[21304]=57;
sine[21305]=57;
sine[21306]=57;
sine[21307]=57;
sine[21308]=57;
sine[21309]=57;
sine[21310]=57;
sine[21311]=57;
sine[21312]=57;
sine[21313]=57;
sine[21314]=57;
sine[21315]=57;
sine[21316]=57;
sine[21317]=58;
sine[21318]=58;
sine[21319]=58;
sine[21320]=58;
sine[21321]=58;
sine[21322]=58;
sine[21323]=58;
sine[21324]=58;
sine[21325]=58;
sine[21326]=58;
sine[21327]=58;
sine[21328]=58;
sine[21329]=58;
sine[21330]=58;
sine[21331]=58;
sine[21332]=58;
sine[21333]=58;
sine[21334]=58;
sine[21335]=58;
sine[21336]=58;
sine[21337]=58;
sine[21338]=58;
sine[21339]=58;
sine[21340]=58;
sine[21341]=58;
sine[21342]=58;
sine[21343]=58;
sine[21344]=58;
sine[21345]=58;
sine[21346]=58;
sine[21347]=59;
sine[21348]=59;
sine[21349]=59;
sine[21350]=59;
sine[21351]=59;
sine[21352]=59;
sine[21353]=59;
sine[21354]=59;
sine[21355]=59;
sine[21356]=59;
sine[21357]=59;
sine[21358]=59;
sine[21359]=59;
sine[21360]=59;
sine[21361]=59;
sine[21362]=59;
sine[21363]=59;
sine[21364]=59;
sine[21365]=59;
sine[21366]=59;
sine[21367]=59;
sine[21368]=59;
sine[21369]=59;
sine[21370]=59;
sine[21371]=59;
sine[21372]=59;
sine[21373]=59;
sine[21374]=59;
sine[21375]=59;
sine[21376]=59;
sine[21377]=59;
sine[21378]=60;
sine[21379]=60;
sine[21380]=60;
sine[21381]=60;
sine[21382]=60;
sine[21383]=60;
sine[21384]=60;
sine[21385]=60;
sine[21386]=60;
sine[21387]=60;
sine[21388]=60;
sine[21389]=60;
sine[21390]=60;
sine[21391]=60;
sine[21392]=60;
sine[21393]=60;
sine[21394]=60;
sine[21395]=60;
sine[21396]=60;
sine[21397]=60;
sine[21398]=60;
sine[21399]=60;
sine[21400]=60;
sine[21401]=60;
sine[21402]=60;
sine[21403]=60;
sine[21404]=60;
sine[21405]=60;
sine[21406]=60;
sine[21407]=60;
sine[21408]=60;
sine[21409]=60;
sine[21410]=61;
sine[21411]=61;
sine[21412]=61;
sine[21413]=61;
sine[21414]=61;
sine[21415]=61;
sine[21416]=61;
sine[21417]=61;
sine[21418]=61;
sine[21419]=61;
sine[21420]=61;
sine[21421]=61;
sine[21422]=61;
sine[21423]=61;
sine[21424]=61;
sine[21425]=61;
sine[21426]=61;
sine[21427]=61;
sine[21428]=61;
sine[21429]=61;
sine[21430]=61;
sine[21431]=61;
sine[21432]=61;
sine[21433]=61;
sine[21434]=61;
sine[21435]=61;
sine[21436]=61;
sine[21437]=61;
sine[21438]=61;
sine[21439]=61;
sine[21440]=61;
sine[21441]=61;
sine[21442]=61;
sine[21443]=62;
sine[21444]=62;
sine[21445]=62;
sine[21446]=62;
sine[21447]=62;
sine[21448]=62;
sine[21449]=62;
sine[21450]=62;
sine[21451]=62;
sine[21452]=62;
sine[21453]=62;
sine[21454]=62;
sine[21455]=62;
sine[21456]=62;
sine[21457]=62;
sine[21458]=62;
sine[21459]=62;
sine[21460]=62;
sine[21461]=62;
sine[21462]=62;
sine[21463]=62;
sine[21464]=62;
sine[21465]=62;
sine[21466]=62;
sine[21467]=62;
sine[21468]=62;
sine[21469]=62;
sine[21470]=62;
sine[21471]=62;
sine[21472]=62;
sine[21473]=62;
sine[21474]=62;
sine[21475]=62;
sine[21476]=63;
sine[21477]=63;
sine[21478]=63;
sine[21479]=63;
sine[21480]=63;
sine[21481]=63;
sine[21482]=63;
sine[21483]=63;
sine[21484]=63;
sine[21485]=63;
sine[21486]=63;
sine[21487]=63;
sine[21488]=63;
sine[21489]=63;
sine[21490]=63;
sine[21491]=63;
sine[21492]=63;
sine[21493]=63;
sine[21494]=63;
sine[21495]=63;
sine[21496]=63;
sine[21497]=63;
sine[21498]=63;
sine[21499]=63;
sine[21500]=63;
sine[21501]=63;
sine[21502]=63;
sine[21503]=63;
sine[21504]=63;
sine[21505]=63;
sine[21506]=63;
sine[21507]=63;
sine[21508]=63;
sine[21509]=63;
sine[21510]=63;
sine[21511]=64;
sine[21512]=64;
sine[21513]=64;
sine[21514]=64;
sine[21515]=64;
sine[21516]=64;
sine[21517]=64;
sine[21518]=64;
sine[21519]=64;
sine[21520]=64;
sine[21521]=64;
sine[21522]=64;
sine[21523]=64;
sine[21524]=64;
sine[21525]=64;
sine[21526]=64;
sine[21527]=64;
sine[21528]=64;
sine[21529]=64;
sine[21530]=64;
sine[21531]=64;
sine[21532]=64;
sine[21533]=64;
sine[21534]=64;
sine[21535]=64;
sine[21536]=64;
sine[21537]=64;
sine[21538]=64;
sine[21539]=64;
sine[21540]=64;
sine[21541]=64;
sine[21542]=64;
sine[21543]=64;
sine[21544]=64;
sine[21545]=64;
sine[21546]=65;
sine[21547]=65;
sine[21548]=65;
sine[21549]=65;
sine[21550]=65;
sine[21551]=65;
sine[21552]=65;
sine[21553]=65;
sine[21554]=65;
sine[21555]=65;
sine[21556]=65;
sine[21557]=65;
sine[21558]=65;
sine[21559]=65;
sine[21560]=65;
sine[21561]=65;
sine[21562]=65;
sine[21563]=65;
sine[21564]=65;
sine[21565]=65;
sine[21566]=65;
sine[21567]=65;
sine[21568]=65;
sine[21569]=65;
sine[21570]=65;
sine[21571]=65;
sine[21572]=65;
sine[21573]=65;
sine[21574]=65;
sine[21575]=65;
sine[21576]=65;
sine[21577]=65;
sine[21578]=65;
sine[21579]=65;
sine[21580]=65;
sine[21581]=65;
sine[21582]=65;
sine[21583]=66;
sine[21584]=66;
sine[21585]=66;
sine[21586]=66;
sine[21587]=66;
sine[21588]=66;
sine[21589]=66;
sine[21590]=66;
sine[21591]=66;
sine[21592]=66;
sine[21593]=66;
sine[21594]=66;
sine[21595]=66;
sine[21596]=66;
sine[21597]=66;
sine[21598]=66;
sine[21599]=66;
sine[21600]=66;
sine[21601]=66;
sine[21602]=66;
sine[21603]=66;
sine[21604]=66;
sine[21605]=66;
sine[21606]=66;
sine[21607]=66;
sine[21608]=66;
sine[21609]=66;
sine[21610]=66;
sine[21611]=66;
sine[21612]=66;
sine[21613]=66;
sine[21614]=66;
sine[21615]=66;
sine[21616]=66;
sine[21617]=66;
sine[21618]=66;
sine[21619]=66;
sine[21620]=66;
sine[21621]=67;
sine[21622]=67;
sine[21623]=67;
sine[21624]=67;
sine[21625]=67;
sine[21626]=67;
sine[21627]=67;
sine[21628]=67;
sine[21629]=67;
sine[21630]=67;
sine[21631]=67;
sine[21632]=67;
sine[21633]=67;
sine[21634]=67;
sine[21635]=67;
sine[21636]=67;
sine[21637]=67;
sine[21638]=67;
sine[21639]=67;
sine[21640]=67;
sine[21641]=67;
sine[21642]=67;
sine[21643]=67;
sine[21644]=67;
sine[21645]=67;
sine[21646]=67;
sine[21647]=67;
sine[21648]=67;
sine[21649]=67;
sine[21650]=67;
sine[21651]=67;
sine[21652]=67;
sine[21653]=67;
sine[21654]=67;
sine[21655]=67;
sine[21656]=67;
sine[21657]=67;
sine[21658]=67;
sine[21659]=67;
sine[21660]=67;
sine[21661]=68;
sine[21662]=68;
sine[21663]=68;
sine[21664]=68;
sine[21665]=68;
sine[21666]=68;
sine[21667]=68;
sine[21668]=68;
sine[21669]=68;
sine[21670]=68;
sine[21671]=68;
sine[21672]=68;
sine[21673]=68;
sine[21674]=68;
sine[21675]=68;
sine[21676]=68;
sine[21677]=68;
sine[21678]=68;
sine[21679]=68;
sine[21680]=68;
sine[21681]=68;
sine[21682]=68;
sine[21683]=68;
sine[21684]=68;
sine[21685]=68;
sine[21686]=68;
sine[21687]=68;
sine[21688]=68;
sine[21689]=68;
sine[21690]=68;
sine[21691]=68;
sine[21692]=68;
sine[21693]=68;
sine[21694]=68;
sine[21695]=68;
sine[21696]=68;
sine[21697]=68;
sine[21698]=68;
sine[21699]=68;
sine[21700]=68;
sine[21701]=68;
sine[21702]=69;
sine[21703]=69;
sine[21704]=69;
sine[21705]=69;
sine[21706]=69;
sine[21707]=69;
sine[21708]=69;
sine[21709]=69;
sine[21710]=69;
sine[21711]=69;
sine[21712]=69;
sine[21713]=69;
sine[21714]=69;
sine[21715]=69;
sine[21716]=69;
sine[21717]=69;
sine[21718]=69;
sine[21719]=69;
sine[21720]=69;
sine[21721]=69;
sine[21722]=69;
sine[21723]=69;
sine[21724]=69;
sine[21725]=69;
sine[21726]=69;
sine[21727]=69;
sine[21728]=69;
sine[21729]=69;
sine[21730]=69;
sine[21731]=69;
sine[21732]=69;
sine[21733]=69;
sine[21734]=69;
sine[21735]=69;
sine[21736]=69;
sine[21737]=69;
sine[21738]=69;
sine[21739]=69;
sine[21740]=69;
sine[21741]=69;
sine[21742]=69;
sine[21743]=69;
sine[21744]=69;
sine[21745]=69;
sine[21746]=70;
sine[21747]=70;
sine[21748]=70;
sine[21749]=70;
sine[21750]=70;
sine[21751]=70;
sine[21752]=70;
sine[21753]=70;
sine[21754]=70;
sine[21755]=70;
sine[21756]=70;
sine[21757]=70;
sine[21758]=70;
sine[21759]=70;
sine[21760]=70;
sine[21761]=70;
sine[21762]=70;
sine[21763]=70;
sine[21764]=70;
sine[21765]=70;
sine[21766]=70;
sine[21767]=70;
sine[21768]=70;
sine[21769]=70;
sine[21770]=70;
sine[21771]=70;
sine[21772]=70;
sine[21773]=70;
sine[21774]=70;
sine[21775]=70;
sine[21776]=70;
sine[21777]=70;
sine[21778]=70;
sine[21779]=70;
sine[21780]=70;
sine[21781]=70;
sine[21782]=70;
sine[21783]=70;
sine[21784]=70;
sine[21785]=70;
sine[21786]=70;
sine[21787]=70;
sine[21788]=70;
sine[21789]=70;
sine[21790]=70;
sine[21791]=71;
sine[21792]=71;
sine[21793]=71;
sine[21794]=71;
sine[21795]=71;
sine[21796]=71;
sine[21797]=71;
sine[21798]=71;
sine[21799]=71;
sine[21800]=71;
sine[21801]=71;
sine[21802]=71;
sine[21803]=71;
sine[21804]=71;
sine[21805]=71;
sine[21806]=71;
sine[21807]=71;
sine[21808]=71;
sine[21809]=71;
sine[21810]=71;
sine[21811]=71;
sine[21812]=71;
sine[21813]=71;
sine[21814]=71;
sine[21815]=71;
sine[21816]=71;
sine[21817]=71;
sine[21818]=71;
sine[21819]=71;
sine[21820]=71;
sine[21821]=71;
sine[21822]=71;
sine[21823]=71;
sine[21824]=71;
sine[21825]=71;
sine[21826]=71;
sine[21827]=71;
sine[21828]=71;
sine[21829]=71;
sine[21830]=71;
sine[21831]=71;
sine[21832]=71;
sine[21833]=71;
sine[21834]=71;
sine[21835]=71;
sine[21836]=71;
sine[21837]=71;
sine[21838]=71;
sine[21839]=71;
sine[21840]=72;
sine[21841]=72;
sine[21842]=72;
sine[21843]=72;
sine[21844]=72;
sine[21845]=72;
sine[21846]=72;
sine[21847]=72;
sine[21848]=72;
sine[21849]=72;
sine[21850]=72;
sine[21851]=72;
sine[21852]=72;
sine[21853]=72;
sine[21854]=72;
sine[21855]=72;
sine[21856]=72;
sine[21857]=72;
sine[21858]=72;
sine[21859]=72;
sine[21860]=72;
sine[21861]=72;
sine[21862]=72;
sine[21863]=72;
sine[21864]=72;
sine[21865]=72;
sine[21866]=72;
sine[21867]=72;
sine[21868]=72;
sine[21869]=72;
sine[21870]=72;
sine[21871]=72;
sine[21872]=72;
sine[21873]=72;
sine[21874]=72;
sine[21875]=72;
sine[21876]=72;
sine[21877]=72;
sine[21878]=72;
sine[21879]=72;
sine[21880]=72;
sine[21881]=72;
sine[21882]=72;
sine[21883]=72;
sine[21884]=72;
sine[21885]=72;
sine[21886]=72;
sine[21887]=72;
sine[21888]=72;
sine[21889]=72;
sine[21890]=72;
sine[21891]=72;
sine[21892]=72;
sine[21893]=73;
sine[21894]=73;
sine[21895]=73;
sine[21896]=73;
sine[21897]=73;
sine[21898]=73;
sine[21899]=73;
sine[21900]=73;
sine[21901]=73;
sine[21902]=73;
sine[21903]=73;
sine[21904]=73;
sine[21905]=73;
sine[21906]=73;
sine[21907]=73;
sine[21908]=73;
sine[21909]=73;
sine[21910]=73;
sine[21911]=73;
sine[21912]=73;
sine[21913]=73;
sine[21914]=73;
sine[21915]=73;
sine[21916]=73;
sine[21917]=73;
sine[21918]=73;
sine[21919]=73;
sine[21920]=73;
sine[21921]=73;
sine[21922]=73;
sine[21923]=73;
sine[21924]=73;
sine[21925]=73;
sine[21926]=73;
sine[21927]=73;
sine[21928]=73;
sine[21929]=73;
sine[21930]=73;
sine[21931]=73;
sine[21932]=73;
sine[21933]=73;
sine[21934]=73;
sine[21935]=73;
sine[21936]=73;
sine[21937]=73;
sine[21938]=73;
sine[21939]=73;
sine[21940]=73;
sine[21941]=73;
sine[21942]=73;
sine[21943]=73;
sine[21944]=73;
sine[21945]=73;
sine[21946]=73;
sine[21947]=73;
sine[21948]=73;
sine[21949]=73;
sine[21950]=74;
sine[21951]=74;
sine[21952]=74;
sine[21953]=74;
sine[21954]=74;
sine[21955]=74;
sine[21956]=74;
sine[21957]=74;
sine[21958]=74;
sine[21959]=74;
sine[21960]=74;
sine[21961]=74;
sine[21962]=74;
sine[21963]=74;
sine[21964]=74;
sine[21965]=74;
sine[21966]=74;
sine[21967]=74;
sine[21968]=74;
sine[21969]=74;
sine[21970]=74;
sine[21971]=74;
sine[21972]=74;
sine[21973]=74;
sine[21974]=74;
sine[21975]=74;
sine[21976]=74;
sine[21977]=74;
sine[21978]=74;
sine[21979]=74;
sine[21980]=74;
sine[21981]=74;
sine[21982]=74;
sine[21983]=74;
sine[21984]=74;
sine[21985]=74;
sine[21986]=74;
sine[21987]=74;
sine[21988]=74;
sine[21989]=74;
sine[21990]=74;
sine[21991]=74;
sine[21992]=74;
sine[21993]=74;
sine[21994]=74;
sine[21995]=74;
sine[21996]=74;
sine[21997]=74;
sine[21998]=74;
sine[21999]=74;
sine[22000]=74;
sine[22001]=74;
sine[22002]=74;
sine[22003]=74;
sine[22004]=74;
sine[22005]=74;
sine[22006]=74;
sine[22007]=74;
sine[22008]=74;
sine[22009]=74;
sine[22010]=74;
sine[22011]=74;
sine[22012]=74;
sine[22013]=74;
sine[22014]=75;
sine[22015]=75;
sine[22016]=75;
sine[22017]=75;
sine[22018]=75;
sine[22019]=75;
sine[22020]=75;
sine[22021]=75;
sine[22022]=75;
sine[22023]=75;
sine[22024]=75;
sine[22025]=75;
sine[22026]=75;
sine[22027]=75;
sine[22028]=75;
sine[22029]=75;
sine[22030]=75;
sine[22031]=75;
sine[22032]=75;
sine[22033]=75;
sine[22034]=75;
sine[22035]=75;
sine[22036]=75;
sine[22037]=75;
sine[22038]=75;
sine[22039]=75;
sine[22040]=75;
sine[22041]=75;
sine[22042]=75;
sine[22043]=75;
sine[22044]=75;
sine[22045]=75;
sine[22046]=75;
sine[22047]=75;
sine[22048]=75;
sine[22049]=75;
sine[22050]=75;
sine[22051]=75;
sine[22052]=75;
sine[22053]=75;
sine[22054]=75;
sine[22055]=75;
sine[22056]=75;
sine[22057]=75;
sine[22058]=75;
sine[22059]=75;
sine[22060]=75;
sine[22061]=75;
sine[22062]=75;
sine[22063]=75;
sine[22064]=75;
sine[22065]=75;
sine[22066]=75;
sine[22067]=75;
sine[22068]=75;
sine[22069]=75;
sine[22070]=75;
sine[22071]=75;
sine[22072]=75;
sine[22073]=75;
sine[22074]=75;
sine[22075]=75;
sine[22076]=75;
sine[22077]=75;
sine[22078]=75;
sine[22079]=75;
sine[22080]=75;
sine[22081]=75;
sine[22082]=75;
sine[22083]=75;
sine[22084]=75;
sine[22085]=75;
sine[22086]=75;
sine[22087]=76;
sine[22088]=76;
sine[22089]=76;
sine[22090]=76;
sine[22091]=76;
sine[22092]=76;
sine[22093]=76;
sine[22094]=76;
sine[22095]=76;
sine[22096]=76;
sine[22097]=76;
sine[22098]=76;
sine[22099]=76;
sine[22100]=76;
sine[22101]=76;
sine[22102]=76;
sine[22103]=76;
sine[22104]=76;
sine[22105]=76;
sine[22106]=76;
sine[22107]=76;
sine[22108]=76;
sine[22109]=76;
sine[22110]=76;
sine[22111]=76;
sine[22112]=76;
sine[22113]=76;
sine[22114]=76;
sine[22115]=76;
sine[22116]=76;
sine[22117]=76;
sine[22118]=76;
sine[22119]=76;
sine[22120]=76;
sine[22121]=76;
sine[22122]=76;
sine[22123]=76;
sine[22124]=76;
sine[22125]=76;
sine[22126]=76;
sine[22127]=76;
sine[22128]=76;
sine[22129]=76;
sine[22130]=76;
sine[22131]=76;
sine[22132]=76;
sine[22133]=76;
sine[22134]=76;
sine[22135]=76;
sine[22136]=76;
sine[22137]=76;
sine[22138]=76;
sine[22139]=76;
sine[22140]=76;
sine[22141]=76;
sine[22142]=76;
sine[22143]=76;
sine[22144]=76;
sine[22145]=76;
sine[22146]=76;
sine[22147]=76;
sine[22148]=76;
sine[22149]=76;
sine[22150]=76;
sine[22151]=76;
sine[22152]=76;
sine[22153]=76;
sine[22154]=76;
sine[22155]=76;
sine[22156]=76;
sine[22157]=76;
sine[22158]=76;
sine[22159]=76;
sine[22160]=76;
sine[22161]=76;
sine[22162]=76;
sine[22163]=76;
sine[22164]=76;
sine[22165]=76;
sine[22166]=76;
sine[22167]=76;
sine[22168]=76;
sine[22169]=76;
sine[22170]=76;
sine[22171]=76;
sine[22172]=76;
sine[22173]=76;
sine[22174]=76;
sine[22175]=77;
sine[22176]=77;
sine[22177]=77;
sine[22178]=77;
sine[22179]=77;
sine[22180]=77;
sine[22181]=77;
sine[22182]=77;
sine[22183]=77;
sine[22184]=77;
sine[22185]=77;
sine[22186]=77;
sine[22187]=77;
sine[22188]=77;
sine[22189]=77;
sine[22190]=77;
sine[22191]=77;
sine[22192]=77;
sine[22193]=77;
sine[22194]=77;
sine[22195]=77;
sine[22196]=77;
sine[22197]=77;
sine[22198]=77;
sine[22199]=77;
sine[22200]=77;
sine[22201]=77;
sine[22202]=77;
sine[22203]=77;
sine[22204]=77;
sine[22205]=77;
sine[22206]=77;
sine[22207]=77;
sine[22208]=77;
sine[22209]=77;
sine[22210]=77;
sine[22211]=77;
sine[22212]=77;
sine[22213]=77;
sine[22214]=77;
sine[22215]=77;
sine[22216]=77;
sine[22217]=77;
sine[22218]=77;
sine[22219]=77;
sine[22220]=77;
sine[22221]=77;
sine[22222]=77;
sine[22223]=77;
sine[22224]=77;
sine[22225]=77;
sine[22226]=77;
sine[22227]=77;
sine[22228]=77;
sine[22229]=77;
sine[22230]=77;
sine[22231]=77;
sine[22232]=77;
sine[22233]=77;
sine[22234]=77;
sine[22235]=77;
sine[22236]=77;
sine[22237]=77;
sine[22238]=77;
sine[22239]=77;
sine[22240]=77;
sine[22241]=77;
sine[22242]=77;
sine[22243]=77;
sine[22244]=77;
sine[22245]=77;
sine[22246]=77;
sine[22247]=77;
sine[22248]=77;
sine[22249]=77;
sine[22250]=77;
sine[22251]=77;
sine[22252]=77;
sine[22253]=77;
sine[22254]=77;
sine[22255]=77;
sine[22256]=77;
sine[22257]=77;
sine[22258]=77;
sine[22259]=77;
sine[22260]=77;
sine[22261]=77;
sine[22262]=77;
sine[22263]=77;
sine[22264]=77;
sine[22265]=77;
sine[22266]=77;
sine[22267]=77;
sine[22268]=77;
sine[22269]=77;
sine[22270]=77;
sine[22271]=77;
sine[22272]=77;
sine[22273]=77;
sine[22274]=77;
sine[22275]=77;
sine[22276]=77;
sine[22277]=77;
sine[22278]=77;
sine[22279]=77;
sine[22280]=77;
sine[22281]=77;
sine[22282]=77;
sine[22283]=77;
sine[22284]=77;
sine[22285]=77;
sine[22286]=77;
sine[22287]=77;
sine[22288]=77;
sine[22289]=77;
sine[22290]=77;
sine[22291]=77;
sine[22292]=77;
sine[22293]=77;
sine[22294]=77;
sine[22295]=77;
sine[22296]=77;
sine[22297]=77;
sine[22298]=77;
sine[22299]=78;
sine[22300]=78;
sine[22301]=78;
sine[22302]=78;
sine[22303]=78;
sine[22304]=78;
sine[22305]=78;
sine[22306]=78;
sine[22307]=78;
sine[22308]=78;
sine[22309]=78;
sine[22310]=78;
sine[22311]=78;
sine[22312]=78;
sine[22313]=78;
sine[22314]=78;
sine[22315]=78;
sine[22316]=78;
sine[22317]=78;
sine[22318]=78;
sine[22319]=78;
sine[22320]=78;
sine[22321]=78;
sine[22322]=78;
sine[22323]=78;
sine[22324]=78;
sine[22325]=78;
sine[22326]=78;
sine[22327]=78;
sine[22328]=78;
sine[22329]=78;
sine[22330]=78;
sine[22331]=78;
sine[22332]=78;
sine[22333]=78;
sine[22334]=78;
sine[22335]=78;
sine[22336]=78;
sine[22337]=78;
sine[22338]=78;
sine[22339]=78;
sine[22340]=78;
sine[22341]=78;
sine[22342]=78;
sine[22343]=78;
sine[22344]=78;
sine[22345]=78;
sine[22346]=78;
sine[22347]=78;
sine[22348]=78;
sine[22349]=78;
sine[22350]=78;
sine[22351]=78;
sine[22352]=78;
sine[22353]=78;
sine[22354]=78;
sine[22355]=78;
sine[22356]=78;
sine[22357]=78;
sine[22358]=78;
sine[22359]=78;
sine[22360]=78;
sine[22361]=78;
sine[22362]=78;
sine[22363]=78;
sine[22364]=78;
sine[22365]=78;
sine[22366]=78;
sine[22367]=78;
sine[22368]=78;
sine[22369]=78;
sine[22370]=78;
sine[22371]=78;
sine[22372]=78;
sine[22373]=78;
sine[22374]=78;
sine[22375]=78;
sine[22376]=78;
sine[22377]=78;
sine[22378]=78;
sine[22379]=78;
sine[22380]=78;
sine[22381]=78;
sine[22382]=78;
sine[22383]=78;
sine[22384]=78;
sine[22385]=78;
sine[22386]=78;
sine[22387]=78;
sine[22388]=78;
sine[22389]=78;
sine[22390]=78;
sine[22391]=78;
sine[22392]=78;
sine[22393]=78;
sine[22394]=78;
sine[22395]=78;
sine[22396]=78;
sine[22397]=78;
sine[22398]=78;
sine[22399]=78;
sine[22400]=78;
sine[22401]=78;
sine[22402]=78;
sine[22403]=78;
sine[22404]=78;
sine[22405]=78;
sine[22406]=78;
sine[22407]=78;
sine[22408]=78;
sine[22409]=78;
sine[22410]=78;
sine[22411]=78;
sine[22412]=78;
sine[22413]=78;
sine[22414]=78;
sine[22415]=78;
sine[22416]=78;
sine[22417]=78;
sine[22418]=78;
sine[22419]=78;
sine[22420]=78;
sine[22421]=78;
sine[22422]=78;
sine[22423]=78;
sine[22424]=78;
sine[22425]=78;
sine[22426]=78;
sine[22427]=78;
sine[22428]=78;
sine[22429]=78;
sine[22430]=78;
sine[22431]=78;
sine[22432]=78;
sine[22433]=78;
sine[22434]=78;
sine[22435]=78;
sine[22436]=78;
sine[22437]=78;
sine[22438]=78;
sine[22439]=78;
sine[22440]=78;
sine[22441]=78;
sine[22442]=78;
sine[22443]=78;
sine[22444]=78;
sine[22445]=78;
sine[22446]=78;
sine[22447]=78;
sine[22448]=78;
sine[22449]=78;
sine[22450]=78;
sine[22451]=78;
sine[22452]=78;
sine[22453]=78;
sine[22454]=78;
sine[22455]=78;
sine[22456]=78;
sine[22457]=78;
sine[22458]=78;
sine[22459]=78;
sine[22460]=78;
sine[22461]=78;
sine[22462]=78;
sine[22463]=78;
sine[22464]=78;
sine[22465]=78;
sine[22466]=78;
sine[22467]=78;
sine[22468]=78;
sine[22469]=78;
sine[22470]=78;
sine[22471]=78;
sine[22472]=78;
sine[22473]=78;
sine[22474]=78;
sine[22475]=78;
sine[22476]=78;
sine[22477]=78;
sine[22478]=78;
sine[22479]=78;
sine[22480]=78;
sine[22481]=78;
sine[22482]=78;
sine[22483]=78;
sine[22484]=78;
sine[22485]=78;
sine[22486]=78;
sine[22487]=78;
sine[22488]=78;
sine[22489]=78;
sine[22490]=78;
sine[22491]=78;
sine[22492]=78;
sine[22493]=78;
sine[22494]=78;
sine[22495]=78;
sine[22496]=78;
sine[22497]=78;
sine[22498]=78;
sine[22499]=78;
sine[22500]=78;
sine[22501]=78;
sine[22502]=78;
sine[22503]=78;
sine[22504]=78;
sine[22505]=78;
sine[22506]=78;
sine[22507]=78;
sine[22508]=78;
sine[22509]=78;
sine[22510]=78;
sine[22511]=78;
sine[22512]=78;
sine[22513]=78;
sine[22514]=78;
sine[22515]=78;
sine[22516]=78;
sine[22517]=78;
sine[22518]=78;
sine[22519]=78;
sine[22520]=78;
sine[22521]=78;
sine[22522]=78;
sine[22523]=78;
sine[22524]=78;
sine[22525]=78;
sine[22526]=78;
sine[22527]=78;
sine[22528]=78;
sine[22529]=78;
sine[22530]=78;
sine[22531]=78;
sine[22532]=78;
sine[22533]=78;
sine[22534]=78;
sine[22535]=78;
sine[22536]=78;
sine[22537]=78;
sine[22538]=78;
sine[22539]=78;
sine[22540]=78;
sine[22541]=78;
sine[22542]=78;
sine[22543]=78;
sine[22544]=78;
sine[22545]=78;
sine[22546]=78;
sine[22547]=78;
sine[22548]=78;
sine[22549]=78;
sine[22550]=78;
sine[22551]=78;
sine[22552]=78;
sine[22553]=78;
sine[22554]=78;
sine[22555]=78;
sine[22556]=78;
sine[22557]=78;
sine[22558]=78;
sine[22559]=78;
sine[22560]=78;
sine[22561]=78;
sine[22562]=78;
sine[22563]=78;
sine[22564]=78;
sine[22565]=78;
sine[22566]=78;
sine[22567]=78;
sine[22568]=78;
sine[22569]=78;
sine[22570]=78;
sine[22571]=78;
sine[22572]=78;
sine[22573]=78;
sine[22574]=78;
sine[22575]=78;
sine[22576]=78;
sine[22577]=78;
sine[22578]=78;
sine[22579]=78;
sine[22580]=78;
sine[22581]=78;
sine[22582]=78;
sine[22583]=78;
sine[22584]=78;
sine[22585]=78;
sine[22586]=78;
sine[22587]=78;
sine[22588]=78;
sine[22589]=78;
sine[22590]=78;
sine[22591]=78;
sine[22592]=78;
sine[22593]=78;
sine[22594]=78;
sine[22595]=78;
sine[22596]=78;
sine[22597]=78;
sine[22598]=78;
sine[22599]=78;
sine[22600]=78;
sine[22601]=78;
sine[22602]=78;
sine[22603]=78;
sine[22604]=78;
sine[22605]=78;
sine[22606]=78;
sine[22607]=78;
sine[22608]=78;
sine[22609]=78;
sine[22610]=78;
sine[22611]=78;
sine[22612]=78;
sine[22613]=78;
sine[22614]=78;
sine[22615]=78;
sine[22616]=78;
sine[22617]=78;
sine[22618]=78;
sine[22619]=78;
sine[22620]=78;
sine[22621]=78;
sine[22622]=78;
sine[22623]=78;
sine[22624]=78;
sine[22625]=78;
sine[22626]=78;
sine[22627]=78;
sine[22628]=78;
sine[22629]=78;
sine[22630]=78;
sine[22631]=78;
sine[22632]=78;
sine[22633]=78;
sine[22634]=78;
sine[22635]=78;
sine[22636]=78;
sine[22637]=78;
sine[22638]=78;
sine[22639]=78;
sine[22640]=78;
sine[22641]=78;
sine[22642]=78;
sine[22643]=78;
sine[22644]=78;
sine[22645]=78;
sine[22646]=78;
sine[22647]=78;
sine[22648]=78;
sine[22649]=78;
sine[22650]=78;
sine[22651]=78;
sine[22652]=78;
sine[22653]=78;
sine[22654]=78;
sine[22655]=78;
sine[22656]=78;
sine[22657]=78;
sine[22658]=78;
sine[22659]=78;
sine[22660]=78;
sine[22661]=78;
sine[22662]=78;
sine[22663]=78;
sine[22664]=78;
sine[22665]=78;
sine[22666]=78;
sine[22667]=78;
sine[22668]=78;
sine[22669]=78;
sine[22670]=78;
sine[22671]=78;
sine[22672]=78;
sine[22673]=78;
sine[22674]=78;
sine[22675]=78;
sine[22676]=78;
sine[22677]=78;
sine[22678]=78;
sine[22679]=78;
sine[22680]=78;
sine[22681]=78;
sine[22682]=78;
sine[22683]=78;
sine[22684]=78;
sine[22685]=78;
sine[22686]=78;
sine[22687]=78;
sine[22688]=78;
sine[22689]=78;
sine[22690]=78;
sine[22691]=78;
sine[22692]=78;
sine[22693]=78;
sine[22694]=78;
sine[22695]=78;
sine[22696]=78;
sine[22697]=78;
sine[22698]=78;
sine[22699]=78;
sine[22700]=78;
sine[22701]=78;
sine[22702]=77;
sine[22703]=77;
sine[22704]=77;
sine[22705]=77;
sine[22706]=77;
sine[22707]=77;
sine[22708]=77;
sine[22709]=77;
sine[22710]=77;
sine[22711]=77;
sine[22712]=77;
sine[22713]=77;
sine[22714]=77;
sine[22715]=77;
sine[22716]=77;
sine[22717]=77;
sine[22718]=77;
sine[22719]=77;
sine[22720]=77;
sine[22721]=77;
sine[22722]=77;
sine[22723]=77;
sine[22724]=77;
sine[22725]=77;
sine[22726]=77;
sine[22727]=77;
sine[22728]=77;
sine[22729]=77;
sine[22730]=77;
sine[22731]=77;
sine[22732]=77;
sine[22733]=77;
sine[22734]=77;
sine[22735]=77;
sine[22736]=77;
sine[22737]=77;
sine[22738]=77;
sine[22739]=77;
sine[22740]=77;
sine[22741]=77;
sine[22742]=77;
sine[22743]=77;
sine[22744]=77;
sine[22745]=77;
sine[22746]=77;
sine[22747]=77;
sine[22748]=77;
sine[22749]=77;
sine[22750]=77;
sine[22751]=77;
sine[22752]=77;
sine[22753]=77;
sine[22754]=77;
sine[22755]=77;
sine[22756]=77;
sine[22757]=77;
sine[22758]=77;
sine[22759]=77;
sine[22760]=77;
sine[22761]=77;
sine[22762]=77;
sine[22763]=77;
sine[22764]=77;
sine[22765]=77;
sine[22766]=77;
sine[22767]=77;
sine[22768]=77;
sine[22769]=77;
sine[22770]=77;
sine[22771]=77;
sine[22772]=77;
sine[22773]=77;
sine[22774]=77;
sine[22775]=77;
sine[22776]=77;
sine[22777]=77;
sine[22778]=77;
sine[22779]=77;
sine[22780]=77;
sine[22781]=77;
sine[22782]=77;
sine[22783]=77;
sine[22784]=77;
sine[22785]=77;
sine[22786]=77;
sine[22787]=77;
sine[22788]=77;
sine[22789]=77;
sine[22790]=77;
sine[22791]=77;
sine[22792]=77;
sine[22793]=77;
sine[22794]=77;
sine[22795]=77;
sine[22796]=77;
sine[22797]=77;
sine[22798]=77;
sine[22799]=77;
sine[22800]=77;
sine[22801]=77;
sine[22802]=77;
sine[22803]=77;
sine[22804]=77;
sine[22805]=77;
sine[22806]=77;
sine[22807]=77;
sine[22808]=77;
sine[22809]=77;
sine[22810]=77;
sine[22811]=77;
sine[22812]=77;
sine[22813]=77;
sine[22814]=77;
sine[22815]=77;
sine[22816]=77;
sine[22817]=77;
sine[22818]=77;
sine[22819]=77;
sine[22820]=77;
sine[22821]=77;
sine[22822]=77;
sine[22823]=77;
sine[22824]=77;
sine[22825]=77;
sine[22826]=76;
sine[22827]=76;
sine[22828]=76;
sine[22829]=76;
sine[22830]=76;
sine[22831]=76;
sine[22832]=76;
sine[22833]=76;
sine[22834]=76;
sine[22835]=76;
sine[22836]=76;
sine[22837]=76;
sine[22838]=76;
sine[22839]=76;
sine[22840]=76;
sine[22841]=76;
sine[22842]=76;
sine[22843]=76;
sine[22844]=76;
sine[22845]=76;
sine[22846]=76;
sine[22847]=76;
sine[22848]=76;
sine[22849]=76;
sine[22850]=76;
sine[22851]=76;
sine[22852]=76;
sine[22853]=76;
sine[22854]=76;
sine[22855]=76;
sine[22856]=76;
sine[22857]=76;
sine[22858]=76;
sine[22859]=76;
sine[22860]=76;
sine[22861]=76;
sine[22862]=76;
sine[22863]=76;
sine[22864]=76;
sine[22865]=76;
sine[22866]=76;
sine[22867]=76;
sine[22868]=76;
sine[22869]=76;
sine[22870]=76;
sine[22871]=76;
sine[22872]=76;
sine[22873]=76;
sine[22874]=76;
sine[22875]=76;
sine[22876]=76;
sine[22877]=76;
sine[22878]=76;
sine[22879]=76;
sine[22880]=76;
sine[22881]=76;
sine[22882]=76;
sine[22883]=76;
sine[22884]=76;
sine[22885]=76;
sine[22886]=76;
sine[22887]=76;
sine[22888]=76;
sine[22889]=76;
sine[22890]=76;
sine[22891]=76;
sine[22892]=76;
sine[22893]=76;
sine[22894]=76;
sine[22895]=76;
sine[22896]=76;
sine[22897]=76;
sine[22898]=76;
sine[22899]=76;
sine[22900]=76;
sine[22901]=76;
sine[22902]=76;
sine[22903]=76;
sine[22904]=76;
sine[22905]=76;
sine[22906]=76;
sine[22907]=76;
sine[22908]=76;
sine[22909]=76;
sine[22910]=76;
sine[22911]=76;
sine[22912]=76;
sine[22913]=76;
sine[22914]=75;
sine[22915]=75;
sine[22916]=75;
sine[22917]=75;
sine[22918]=75;
sine[22919]=75;
sine[22920]=75;
sine[22921]=75;
sine[22922]=75;
sine[22923]=75;
sine[22924]=75;
sine[22925]=75;
sine[22926]=75;
sine[22927]=75;
sine[22928]=75;
sine[22929]=75;
sine[22930]=75;
sine[22931]=75;
sine[22932]=75;
sine[22933]=75;
sine[22934]=75;
sine[22935]=75;
sine[22936]=75;
sine[22937]=75;
sine[22938]=75;
sine[22939]=75;
sine[22940]=75;
sine[22941]=75;
sine[22942]=75;
sine[22943]=75;
sine[22944]=75;
sine[22945]=75;
sine[22946]=75;
sine[22947]=75;
sine[22948]=75;
sine[22949]=75;
sine[22950]=75;
sine[22951]=75;
sine[22952]=75;
sine[22953]=75;
sine[22954]=75;
sine[22955]=75;
sine[22956]=75;
sine[22957]=75;
sine[22958]=75;
sine[22959]=75;
sine[22960]=75;
sine[22961]=75;
sine[22962]=75;
sine[22963]=75;
sine[22964]=75;
sine[22965]=75;
sine[22966]=75;
sine[22967]=75;
sine[22968]=75;
sine[22969]=75;
sine[22970]=75;
sine[22971]=75;
sine[22972]=75;
sine[22973]=75;
sine[22974]=75;
sine[22975]=75;
sine[22976]=75;
sine[22977]=75;
sine[22978]=75;
sine[22979]=75;
sine[22980]=75;
sine[22981]=75;
sine[22982]=75;
sine[22983]=75;
sine[22984]=75;
sine[22985]=75;
sine[22986]=75;
sine[22987]=74;
sine[22988]=74;
sine[22989]=74;
sine[22990]=74;
sine[22991]=74;
sine[22992]=74;
sine[22993]=74;
sine[22994]=74;
sine[22995]=74;
sine[22996]=74;
sine[22997]=74;
sine[22998]=74;
sine[22999]=74;
sine[23000]=74;
sine[23001]=74;
sine[23002]=74;
sine[23003]=74;
sine[23004]=74;
sine[23005]=74;
sine[23006]=74;
sine[23007]=74;
sine[23008]=74;
sine[23009]=74;
sine[23010]=74;
sine[23011]=74;
sine[23012]=74;
sine[23013]=74;
sine[23014]=74;
sine[23015]=74;
sine[23016]=74;
sine[23017]=74;
sine[23018]=74;
sine[23019]=74;
sine[23020]=74;
sine[23021]=74;
sine[23022]=74;
sine[23023]=74;
sine[23024]=74;
sine[23025]=74;
sine[23026]=74;
sine[23027]=74;
sine[23028]=74;
sine[23029]=74;
sine[23030]=74;
sine[23031]=74;
sine[23032]=74;
sine[23033]=74;
sine[23034]=74;
sine[23035]=74;
sine[23036]=74;
sine[23037]=74;
sine[23038]=74;
sine[23039]=74;
sine[23040]=74;
sine[23041]=74;
sine[23042]=74;
sine[23043]=74;
sine[23044]=74;
sine[23045]=74;
sine[23046]=74;
sine[23047]=74;
sine[23048]=74;
sine[23049]=74;
sine[23050]=74;
sine[23051]=73;
sine[23052]=73;
sine[23053]=73;
sine[23054]=73;
sine[23055]=73;
sine[23056]=73;
sine[23057]=73;
sine[23058]=73;
sine[23059]=73;
sine[23060]=73;
sine[23061]=73;
sine[23062]=73;
sine[23063]=73;
sine[23064]=73;
sine[23065]=73;
sine[23066]=73;
sine[23067]=73;
sine[23068]=73;
sine[23069]=73;
sine[23070]=73;
sine[23071]=73;
sine[23072]=73;
sine[23073]=73;
sine[23074]=73;
sine[23075]=73;
sine[23076]=73;
sine[23077]=73;
sine[23078]=73;
sine[23079]=73;
sine[23080]=73;
sine[23081]=73;
sine[23082]=73;
sine[23083]=73;
sine[23084]=73;
sine[23085]=73;
sine[23086]=73;
sine[23087]=73;
sine[23088]=73;
sine[23089]=73;
sine[23090]=73;
sine[23091]=73;
sine[23092]=73;
sine[23093]=73;
sine[23094]=73;
sine[23095]=73;
sine[23096]=73;
sine[23097]=73;
sine[23098]=73;
sine[23099]=73;
sine[23100]=73;
sine[23101]=73;
sine[23102]=73;
sine[23103]=73;
sine[23104]=73;
sine[23105]=73;
sine[23106]=73;
sine[23107]=73;
sine[23108]=72;
sine[23109]=72;
sine[23110]=72;
sine[23111]=72;
sine[23112]=72;
sine[23113]=72;
sine[23114]=72;
sine[23115]=72;
sine[23116]=72;
sine[23117]=72;
sine[23118]=72;
sine[23119]=72;
sine[23120]=72;
sine[23121]=72;
sine[23122]=72;
sine[23123]=72;
sine[23124]=72;
sine[23125]=72;
sine[23126]=72;
sine[23127]=72;
sine[23128]=72;
sine[23129]=72;
sine[23130]=72;
sine[23131]=72;
sine[23132]=72;
sine[23133]=72;
sine[23134]=72;
sine[23135]=72;
sine[23136]=72;
sine[23137]=72;
sine[23138]=72;
sine[23139]=72;
sine[23140]=72;
sine[23141]=72;
sine[23142]=72;
sine[23143]=72;
sine[23144]=72;
sine[23145]=72;
sine[23146]=72;
sine[23147]=72;
sine[23148]=72;
sine[23149]=72;
sine[23150]=72;
sine[23151]=72;
sine[23152]=72;
sine[23153]=72;
sine[23154]=72;
sine[23155]=72;
sine[23156]=72;
sine[23157]=72;
sine[23158]=72;
sine[23159]=72;
sine[23160]=72;
sine[23161]=71;
sine[23162]=71;
sine[23163]=71;
sine[23164]=71;
sine[23165]=71;
sine[23166]=71;
sine[23167]=71;
sine[23168]=71;
sine[23169]=71;
sine[23170]=71;
sine[23171]=71;
sine[23172]=71;
sine[23173]=71;
sine[23174]=71;
sine[23175]=71;
sine[23176]=71;
sine[23177]=71;
sine[23178]=71;
sine[23179]=71;
sine[23180]=71;
sine[23181]=71;
sine[23182]=71;
sine[23183]=71;
sine[23184]=71;
sine[23185]=71;
sine[23186]=71;
sine[23187]=71;
sine[23188]=71;
sine[23189]=71;
sine[23190]=71;
sine[23191]=71;
sine[23192]=71;
sine[23193]=71;
sine[23194]=71;
sine[23195]=71;
sine[23196]=71;
sine[23197]=71;
sine[23198]=71;
sine[23199]=71;
sine[23200]=71;
sine[23201]=71;
sine[23202]=71;
sine[23203]=71;
sine[23204]=71;
sine[23205]=71;
sine[23206]=71;
sine[23207]=71;
sine[23208]=71;
sine[23209]=71;
sine[23210]=70;
sine[23211]=70;
sine[23212]=70;
sine[23213]=70;
sine[23214]=70;
sine[23215]=70;
sine[23216]=70;
sine[23217]=70;
sine[23218]=70;
sine[23219]=70;
sine[23220]=70;
sine[23221]=70;
sine[23222]=70;
sine[23223]=70;
sine[23224]=70;
sine[23225]=70;
sine[23226]=70;
sine[23227]=70;
sine[23228]=70;
sine[23229]=70;
sine[23230]=70;
sine[23231]=70;
sine[23232]=70;
sine[23233]=70;
sine[23234]=70;
sine[23235]=70;
sine[23236]=70;
sine[23237]=70;
sine[23238]=70;
sine[23239]=70;
sine[23240]=70;
sine[23241]=70;
sine[23242]=70;
sine[23243]=70;
sine[23244]=70;
sine[23245]=70;
sine[23246]=70;
sine[23247]=70;
sine[23248]=70;
sine[23249]=70;
sine[23250]=70;
sine[23251]=70;
sine[23252]=70;
sine[23253]=70;
sine[23254]=70;
sine[23255]=69;
sine[23256]=69;
sine[23257]=69;
sine[23258]=69;
sine[23259]=69;
sine[23260]=69;
sine[23261]=69;
sine[23262]=69;
sine[23263]=69;
sine[23264]=69;
sine[23265]=69;
sine[23266]=69;
sine[23267]=69;
sine[23268]=69;
sine[23269]=69;
sine[23270]=69;
sine[23271]=69;
sine[23272]=69;
sine[23273]=69;
sine[23274]=69;
sine[23275]=69;
sine[23276]=69;
sine[23277]=69;
sine[23278]=69;
sine[23279]=69;
sine[23280]=69;
sine[23281]=69;
sine[23282]=69;
sine[23283]=69;
sine[23284]=69;
sine[23285]=69;
sine[23286]=69;
sine[23287]=69;
sine[23288]=69;
sine[23289]=69;
sine[23290]=69;
sine[23291]=69;
sine[23292]=69;
sine[23293]=69;
sine[23294]=69;
sine[23295]=69;
sine[23296]=69;
sine[23297]=69;
sine[23298]=69;
sine[23299]=68;
sine[23300]=68;
sine[23301]=68;
sine[23302]=68;
sine[23303]=68;
sine[23304]=68;
sine[23305]=68;
sine[23306]=68;
sine[23307]=68;
sine[23308]=68;
sine[23309]=68;
sine[23310]=68;
sine[23311]=68;
sine[23312]=68;
sine[23313]=68;
sine[23314]=68;
sine[23315]=68;
sine[23316]=68;
sine[23317]=68;
sine[23318]=68;
sine[23319]=68;
sine[23320]=68;
sine[23321]=68;
sine[23322]=68;
sine[23323]=68;
sine[23324]=68;
sine[23325]=68;
sine[23326]=68;
sine[23327]=68;
sine[23328]=68;
sine[23329]=68;
sine[23330]=68;
sine[23331]=68;
sine[23332]=68;
sine[23333]=68;
sine[23334]=68;
sine[23335]=68;
sine[23336]=68;
sine[23337]=68;
sine[23338]=68;
sine[23339]=68;
sine[23340]=67;
sine[23341]=67;
sine[23342]=67;
sine[23343]=67;
sine[23344]=67;
sine[23345]=67;
sine[23346]=67;
sine[23347]=67;
sine[23348]=67;
sine[23349]=67;
sine[23350]=67;
sine[23351]=67;
sine[23352]=67;
sine[23353]=67;
sine[23354]=67;
sine[23355]=67;
sine[23356]=67;
sine[23357]=67;
sine[23358]=67;
sine[23359]=67;
sine[23360]=67;
sine[23361]=67;
sine[23362]=67;
sine[23363]=67;
sine[23364]=67;
sine[23365]=67;
sine[23366]=67;
sine[23367]=67;
sine[23368]=67;
sine[23369]=67;
sine[23370]=67;
sine[23371]=67;
sine[23372]=67;
sine[23373]=67;
sine[23374]=67;
sine[23375]=67;
sine[23376]=67;
sine[23377]=67;
sine[23378]=67;
sine[23379]=67;
sine[23380]=66;
sine[23381]=66;
sine[23382]=66;
sine[23383]=66;
sine[23384]=66;
sine[23385]=66;
sine[23386]=66;
sine[23387]=66;
sine[23388]=66;
sine[23389]=66;
sine[23390]=66;
sine[23391]=66;
sine[23392]=66;
sine[23393]=66;
sine[23394]=66;
sine[23395]=66;
sine[23396]=66;
sine[23397]=66;
sine[23398]=66;
sine[23399]=66;
sine[23400]=66;
sine[23401]=66;
sine[23402]=66;
sine[23403]=66;
sine[23404]=66;
sine[23405]=66;
sine[23406]=66;
sine[23407]=66;
sine[23408]=66;
sine[23409]=66;
sine[23410]=66;
sine[23411]=66;
sine[23412]=66;
sine[23413]=66;
sine[23414]=66;
sine[23415]=66;
sine[23416]=66;
sine[23417]=66;
sine[23418]=65;
sine[23419]=65;
sine[23420]=65;
sine[23421]=65;
sine[23422]=65;
sine[23423]=65;
sine[23424]=65;
sine[23425]=65;
sine[23426]=65;
sine[23427]=65;
sine[23428]=65;
sine[23429]=65;
sine[23430]=65;
sine[23431]=65;
sine[23432]=65;
sine[23433]=65;
sine[23434]=65;
sine[23435]=65;
sine[23436]=65;
sine[23437]=65;
sine[23438]=65;
sine[23439]=65;
sine[23440]=65;
sine[23441]=65;
sine[23442]=65;
sine[23443]=65;
sine[23444]=65;
sine[23445]=65;
sine[23446]=65;
sine[23447]=65;
sine[23448]=65;
sine[23449]=65;
sine[23450]=65;
sine[23451]=65;
sine[23452]=65;
sine[23453]=65;
sine[23454]=65;
sine[23455]=64;
sine[23456]=64;
sine[23457]=64;
sine[23458]=64;
sine[23459]=64;
sine[23460]=64;
sine[23461]=64;
sine[23462]=64;
sine[23463]=64;
sine[23464]=64;
sine[23465]=64;
sine[23466]=64;
sine[23467]=64;
sine[23468]=64;
sine[23469]=64;
sine[23470]=64;
sine[23471]=64;
sine[23472]=64;
sine[23473]=64;
sine[23474]=64;
sine[23475]=64;
sine[23476]=64;
sine[23477]=64;
sine[23478]=64;
sine[23479]=64;
sine[23480]=64;
sine[23481]=64;
sine[23482]=64;
sine[23483]=64;
sine[23484]=64;
sine[23485]=64;
sine[23486]=64;
sine[23487]=64;
sine[23488]=64;
sine[23489]=64;
sine[23490]=63;
sine[23491]=63;
sine[23492]=63;
sine[23493]=63;
sine[23494]=63;
sine[23495]=63;
sine[23496]=63;
sine[23497]=63;
sine[23498]=63;
sine[23499]=63;
sine[23500]=63;
sine[23501]=63;
sine[23502]=63;
sine[23503]=63;
sine[23504]=63;
sine[23505]=63;
sine[23506]=63;
sine[23507]=63;
sine[23508]=63;
sine[23509]=63;
sine[23510]=63;
sine[23511]=63;
sine[23512]=63;
sine[23513]=63;
sine[23514]=63;
sine[23515]=63;
sine[23516]=63;
sine[23517]=63;
sine[23518]=63;
sine[23519]=63;
sine[23520]=63;
sine[23521]=63;
sine[23522]=63;
sine[23523]=63;
sine[23524]=63;
sine[23525]=62;
sine[23526]=62;
sine[23527]=62;
sine[23528]=62;
sine[23529]=62;
sine[23530]=62;
sine[23531]=62;
sine[23532]=62;
sine[23533]=62;
sine[23534]=62;
sine[23535]=62;
sine[23536]=62;
sine[23537]=62;
sine[23538]=62;
sine[23539]=62;
sine[23540]=62;
sine[23541]=62;
sine[23542]=62;
sine[23543]=62;
sine[23544]=62;
sine[23545]=62;
sine[23546]=62;
sine[23547]=62;
sine[23548]=62;
sine[23549]=62;
sine[23550]=62;
sine[23551]=62;
sine[23552]=62;
sine[23553]=62;
sine[23554]=62;
sine[23555]=62;
sine[23556]=62;
sine[23557]=62;
sine[23558]=61;
sine[23559]=61;
sine[23560]=61;
sine[23561]=61;
sine[23562]=61;
sine[23563]=61;
sine[23564]=61;
sine[23565]=61;
sine[23566]=61;
sine[23567]=61;
sine[23568]=61;
sine[23569]=61;
sine[23570]=61;
sine[23571]=61;
sine[23572]=61;
sine[23573]=61;
sine[23574]=61;
sine[23575]=61;
sine[23576]=61;
sine[23577]=61;
sine[23578]=61;
sine[23579]=61;
sine[23580]=61;
sine[23581]=61;
sine[23582]=61;
sine[23583]=61;
sine[23584]=61;
sine[23585]=61;
sine[23586]=61;
sine[23587]=61;
sine[23588]=61;
sine[23589]=61;
sine[23590]=61;
sine[23591]=60;
sine[23592]=60;
sine[23593]=60;
sine[23594]=60;
sine[23595]=60;
sine[23596]=60;
sine[23597]=60;
sine[23598]=60;
sine[23599]=60;
sine[23600]=60;
sine[23601]=60;
sine[23602]=60;
sine[23603]=60;
sine[23604]=60;
sine[23605]=60;
sine[23606]=60;
sine[23607]=60;
sine[23608]=60;
sine[23609]=60;
sine[23610]=60;
sine[23611]=60;
sine[23612]=60;
sine[23613]=60;
sine[23614]=60;
sine[23615]=60;
sine[23616]=60;
sine[23617]=60;
sine[23618]=60;
sine[23619]=60;
sine[23620]=60;
sine[23621]=60;
sine[23622]=60;
sine[23623]=59;
sine[23624]=59;
sine[23625]=59;
sine[23626]=59;
sine[23627]=59;
sine[23628]=59;
sine[23629]=59;
sine[23630]=59;
sine[23631]=59;
sine[23632]=59;
sine[23633]=59;
sine[23634]=59;
sine[23635]=59;
sine[23636]=59;
sine[23637]=59;
sine[23638]=59;
sine[23639]=59;
sine[23640]=59;
sine[23641]=59;
sine[23642]=59;
sine[23643]=59;
sine[23644]=59;
sine[23645]=59;
sine[23646]=59;
sine[23647]=59;
sine[23648]=59;
sine[23649]=59;
sine[23650]=59;
sine[23651]=59;
sine[23652]=59;
sine[23653]=59;
sine[23654]=58;
sine[23655]=58;
sine[23656]=58;
sine[23657]=58;
sine[23658]=58;
sine[23659]=58;
sine[23660]=58;
sine[23661]=58;
sine[23662]=58;
sine[23663]=58;
sine[23664]=58;
sine[23665]=58;
sine[23666]=58;
sine[23667]=58;
sine[23668]=58;
sine[23669]=58;
sine[23670]=58;
sine[23671]=58;
sine[23672]=58;
sine[23673]=58;
sine[23674]=58;
sine[23675]=58;
sine[23676]=58;
sine[23677]=58;
sine[23678]=58;
sine[23679]=58;
sine[23680]=58;
sine[23681]=58;
sine[23682]=58;
sine[23683]=58;
sine[23684]=57;
sine[23685]=57;
sine[23686]=57;
sine[23687]=57;
sine[23688]=57;
sine[23689]=57;
sine[23690]=57;
sine[23691]=57;
sine[23692]=57;
sine[23693]=57;
sine[23694]=57;
sine[23695]=57;
sine[23696]=57;
sine[23697]=57;
sine[23698]=57;
sine[23699]=57;
sine[23700]=57;
sine[23701]=57;
sine[23702]=57;
sine[23703]=57;
sine[23704]=57;
sine[23705]=57;
sine[23706]=57;
sine[23707]=57;
sine[23708]=57;
sine[23709]=57;
sine[23710]=57;
sine[23711]=57;
sine[23712]=57;
sine[23713]=57;
sine[23714]=56;
sine[23715]=56;
sine[23716]=56;
sine[23717]=56;
sine[23718]=56;
sine[23719]=56;
sine[23720]=56;
sine[23721]=56;
sine[23722]=56;
sine[23723]=56;
sine[23724]=56;
sine[23725]=56;
sine[23726]=56;
sine[23727]=56;
sine[23728]=56;
sine[23729]=56;
sine[23730]=56;
sine[23731]=56;
sine[23732]=56;
sine[23733]=56;
sine[23734]=56;
sine[23735]=56;
sine[23736]=56;
sine[23737]=56;
sine[23738]=56;
sine[23739]=56;
sine[23740]=56;
sine[23741]=56;
sine[23742]=56;
sine[23743]=55;
sine[23744]=55;
sine[23745]=55;
sine[23746]=55;
sine[23747]=55;
sine[23748]=55;
sine[23749]=55;
sine[23750]=55;
sine[23751]=55;
sine[23752]=55;
sine[23753]=55;
sine[23754]=55;
sine[23755]=55;
sine[23756]=55;
sine[23757]=55;
sine[23758]=55;
sine[23759]=55;
sine[23760]=55;
sine[23761]=55;
sine[23762]=55;
sine[23763]=55;
sine[23764]=55;
sine[23765]=55;
sine[23766]=55;
sine[23767]=55;
sine[23768]=55;
sine[23769]=55;
sine[23770]=55;
sine[23771]=55;
sine[23772]=54;
sine[23773]=54;
sine[23774]=54;
sine[23775]=54;
sine[23776]=54;
sine[23777]=54;
sine[23778]=54;
sine[23779]=54;
sine[23780]=54;
sine[23781]=54;
sine[23782]=54;
sine[23783]=54;
sine[23784]=54;
sine[23785]=54;
sine[23786]=54;
sine[23787]=54;
sine[23788]=54;
sine[23789]=54;
sine[23790]=54;
sine[23791]=54;
sine[23792]=54;
sine[23793]=54;
sine[23794]=54;
sine[23795]=54;
sine[23796]=54;
sine[23797]=54;
sine[23798]=54;
sine[23799]=54;
sine[23800]=53;
sine[23801]=53;
sine[23802]=53;
sine[23803]=53;
sine[23804]=53;
sine[23805]=53;
sine[23806]=53;
sine[23807]=53;
sine[23808]=53;
sine[23809]=53;
sine[23810]=53;
sine[23811]=53;
sine[23812]=53;
sine[23813]=53;
sine[23814]=53;
sine[23815]=53;
sine[23816]=53;
sine[23817]=53;
sine[23818]=53;
sine[23819]=53;
sine[23820]=53;
sine[23821]=53;
sine[23822]=53;
sine[23823]=53;
sine[23824]=53;
sine[23825]=53;
sine[23826]=53;
sine[23827]=53;
sine[23828]=52;
sine[23829]=52;
sine[23830]=52;
sine[23831]=52;
sine[23832]=52;
sine[23833]=52;
sine[23834]=52;
sine[23835]=52;
sine[23836]=52;
sine[23837]=52;
sine[23838]=52;
sine[23839]=52;
sine[23840]=52;
sine[23841]=52;
sine[23842]=52;
sine[23843]=52;
sine[23844]=52;
sine[23845]=52;
sine[23846]=52;
sine[23847]=52;
sine[23848]=52;
sine[23849]=52;
sine[23850]=52;
sine[23851]=52;
sine[23852]=52;
sine[23853]=52;
sine[23854]=52;
sine[23855]=51;
sine[23856]=51;
sine[23857]=51;
sine[23858]=51;
sine[23859]=51;
sine[23860]=51;
sine[23861]=51;
sine[23862]=51;
sine[23863]=51;
sine[23864]=51;
sine[23865]=51;
sine[23866]=51;
sine[23867]=51;
sine[23868]=51;
sine[23869]=51;
sine[23870]=51;
sine[23871]=51;
sine[23872]=51;
sine[23873]=51;
sine[23874]=51;
sine[23875]=51;
sine[23876]=51;
sine[23877]=51;
sine[23878]=51;
sine[23879]=51;
sine[23880]=51;
sine[23881]=51;
sine[23882]=50;
sine[23883]=50;
sine[23884]=50;
sine[23885]=50;
sine[23886]=50;
sine[23887]=50;
sine[23888]=50;
sine[23889]=50;
sine[23890]=50;
sine[23891]=50;
sine[23892]=50;
sine[23893]=50;
sine[23894]=50;
sine[23895]=50;
sine[23896]=50;
sine[23897]=50;
sine[23898]=50;
sine[23899]=50;
sine[23900]=50;
sine[23901]=50;
sine[23902]=50;
sine[23903]=50;
sine[23904]=50;
sine[23905]=50;
sine[23906]=50;
sine[23907]=50;
sine[23908]=49;
sine[23909]=49;
sine[23910]=49;
sine[23911]=49;
sine[23912]=49;
sine[23913]=49;
sine[23914]=49;
sine[23915]=49;
sine[23916]=49;
sine[23917]=49;
sine[23918]=49;
sine[23919]=49;
sine[23920]=49;
sine[23921]=49;
sine[23922]=49;
sine[23923]=49;
sine[23924]=49;
sine[23925]=49;
sine[23926]=49;
sine[23927]=49;
sine[23928]=49;
sine[23929]=49;
sine[23930]=49;
sine[23931]=49;
sine[23932]=49;
sine[23933]=49;
sine[23934]=49;
sine[23935]=48;
sine[23936]=48;
sine[23937]=48;
sine[23938]=48;
sine[23939]=48;
sine[23940]=48;
sine[23941]=48;
sine[23942]=48;
sine[23943]=48;
sine[23944]=48;
sine[23945]=48;
sine[23946]=48;
sine[23947]=48;
sine[23948]=48;
sine[23949]=48;
sine[23950]=48;
sine[23951]=48;
sine[23952]=48;
sine[23953]=48;
sine[23954]=48;
sine[23955]=48;
sine[23956]=48;
sine[23957]=48;
sine[23958]=48;
sine[23959]=48;
sine[23960]=47;
sine[23961]=47;
sine[23962]=47;
sine[23963]=47;
sine[23964]=47;
sine[23965]=47;
sine[23966]=47;
sine[23967]=47;
sine[23968]=47;
sine[23969]=47;
sine[23970]=47;
sine[23971]=47;
sine[23972]=47;
sine[23973]=47;
sine[23974]=47;
sine[23975]=47;
sine[23976]=47;
sine[23977]=47;
sine[23978]=47;
sine[23979]=47;
sine[23980]=47;
sine[23981]=47;
sine[23982]=47;
sine[23983]=47;
sine[23984]=47;
sine[23985]=47;
sine[23986]=46;
sine[23987]=46;
sine[23988]=46;
sine[23989]=46;
sine[23990]=46;
sine[23991]=46;
sine[23992]=46;
sine[23993]=46;
sine[23994]=46;
sine[23995]=46;
sine[23996]=46;
sine[23997]=46;
sine[23998]=46;
sine[23999]=46;
sine[24000]=46;
sine[24001]=46;
sine[24002]=46;
sine[24003]=46;
sine[24004]=46;
sine[24005]=46;
sine[24006]=46;
sine[24007]=46;
sine[24008]=46;
sine[24009]=46;
sine[24010]=46;
sine[24011]=45;
sine[24012]=45;
sine[24013]=45;
sine[24014]=45;
sine[24015]=45;
sine[24016]=45;
sine[24017]=45;
sine[24018]=45;
sine[24019]=45;
sine[24020]=45;
sine[24021]=45;
sine[24022]=45;
sine[24023]=45;
sine[24024]=45;
sine[24025]=45;
sine[24026]=45;
sine[24027]=45;
sine[24028]=45;
sine[24029]=45;
sine[24030]=45;
sine[24031]=45;
sine[24032]=45;
sine[24033]=45;
sine[24034]=45;
sine[24035]=45;
sine[24036]=44;
sine[24037]=44;
sine[24038]=44;
sine[24039]=44;
sine[24040]=44;
sine[24041]=44;
sine[24042]=44;
sine[24043]=44;
sine[24044]=44;
sine[24045]=44;
sine[24046]=44;
sine[24047]=44;
sine[24048]=44;
sine[24049]=44;
sine[24050]=44;
sine[24051]=44;
sine[24052]=44;
sine[24053]=44;
sine[24054]=44;
sine[24055]=44;
sine[24056]=44;
sine[24057]=44;
sine[24058]=44;
sine[24059]=44;
sine[24060]=44;
sine[24061]=43;
sine[24062]=43;
sine[24063]=43;
sine[24064]=43;
sine[24065]=43;
sine[24066]=43;
sine[24067]=43;
sine[24068]=43;
sine[24069]=43;
sine[24070]=43;
sine[24071]=43;
sine[24072]=43;
sine[24073]=43;
sine[24074]=43;
sine[24075]=43;
sine[24076]=43;
sine[24077]=43;
sine[24078]=43;
sine[24079]=43;
sine[24080]=43;
sine[24081]=43;
sine[24082]=43;
sine[24083]=43;
sine[24084]=43;
sine[24085]=42;
sine[24086]=42;
sine[24087]=42;
sine[24088]=42;
sine[24089]=42;
sine[24090]=42;
sine[24091]=42;
sine[24092]=42;
sine[24093]=42;
sine[24094]=42;
sine[24095]=42;
sine[24096]=42;
sine[24097]=42;
sine[24098]=42;
sine[24099]=42;
sine[24100]=42;
sine[24101]=42;
sine[24102]=42;
sine[24103]=42;
sine[24104]=42;
sine[24105]=42;
sine[24106]=42;
sine[24107]=42;
sine[24108]=42;
sine[24109]=41;
sine[24110]=41;
sine[24111]=41;
sine[24112]=41;
sine[24113]=41;
sine[24114]=41;
sine[24115]=41;
sine[24116]=41;
sine[24117]=41;
sine[24118]=41;
sine[24119]=41;
sine[24120]=41;
sine[24121]=41;
sine[24122]=41;
sine[24123]=41;
sine[24124]=41;
sine[24125]=41;
sine[24126]=41;
sine[24127]=41;
sine[24128]=41;
sine[24129]=41;
sine[24130]=41;
sine[24131]=41;
sine[24132]=41;
sine[24133]=40;
sine[24134]=40;
sine[24135]=40;
sine[24136]=40;
sine[24137]=40;
sine[24138]=40;
sine[24139]=40;
sine[24140]=40;
sine[24141]=40;
sine[24142]=40;
sine[24143]=40;
sine[24144]=40;
sine[24145]=40;
sine[24146]=40;
sine[24147]=40;
sine[24148]=40;
sine[24149]=40;
sine[24150]=40;
sine[24151]=40;
sine[24152]=40;
sine[24153]=40;
sine[24154]=40;
sine[24155]=40;
sine[24156]=40;
sine[24157]=39;
sine[24158]=39;
sine[24159]=39;
sine[24160]=39;
sine[24161]=39;
sine[24162]=39;
sine[24163]=39;
sine[24164]=39;
sine[24165]=39;
sine[24166]=39;
sine[24167]=39;
sine[24168]=39;
sine[24169]=39;
sine[24170]=39;
sine[24171]=39;
sine[24172]=39;
sine[24173]=39;
sine[24174]=39;
sine[24175]=39;
sine[24176]=39;
sine[24177]=39;
sine[24178]=39;
sine[24179]=39;
sine[24180]=38;
sine[24181]=38;
sine[24182]=38;
sine[24183]=38;
sine[24184]=38;
sine[24185]=38;
sine[24186]=38;
sine[24187]=38;
sine[24188]=38;
sine[24189]=38;
sine[24190]=38;
sine[24191]=38;
sine[24192]=38;
sine[24193]=38;
sine[24194]=38;
sine[24195]=38;
sine[24196]=38;
sine[24197]=38;
sine[24198]=38;
sine[24199]=38;
sine[24200]=38;
sine[24201]=38;
sine[24202]=38;
sine[24203]=38;
sine[24204]=37;
sine[24205]=37;
sine[24206]=37;
sine[24207]=37;
sine[24208]=37;
sine[24209]=37;
sine[24210]=37;
sine[24211]=37;
sine[24212]=37;
sine[24213]=37;
sine[24214]=37;
sine[24215]=37;
sine[24216]=37;
sine[24217]=37;
sine[24218]=37;
sine[24219]=37;
sine[24220]=37;
sine[24221]=37;
sine[24222]=37;
sine[24223]=37;
sine[24224]=37;
sine[24225]=37;
sine[24226]=37;
sine[24227]=36;
sine[24228]=36;
sine[24229]=36;
sine[24230]=36;
sine[24231]=36;
sine[24232]=36;
sine[24233]=36;
sine[24234]=36;
sine[24235]=36;
sine[24236]=36;
sine[24237]=36;
sine[24238]=36;
sine[24239]=36;
sine[24240]=36;
sine[24241]=36;
sine[24242]=36;
sine[24243]=36;
sine[24244]=36;
sine[24245]=36;
sine[24246]=36;
sine[24247]=36;
sine[24248]=36;
sine[24249]=36;
sine[24250]=35;
sine[24251]=35;
sine[24252]=35;
sine[24253]=35;
sine[24254]=35;
sine[24255]=35;
sine[24256]=35;
sine[24257]=35;
sine[24258]=35;
sine[24259]=35;
sine[24260]=35;
sine[24261]=35;
sine[24262]=35;
sine[24263]=35;
sine[24264]=35;
sine[24265]=35;
sine[24266]=35;
sine[24267]=35;
sine[24268]=35;
sine[24269]=35;
sine[24270]=35;
sine[24271]=35;
sine[24272]=35;
sine[24273]=34;
sine[24274]=34;
sine[24275]=34;
sine[24276]=34;
sine[24277]=34;
sine[24278]=34;
sine[24279]=34;
sine[24280]=34;
sine[24281]=34;
sine[24282]=34;
sine[24283]=34;
sine[24284]=34;
sine[24285]=34;
sine[24286]=34;
sine[24287]=34;
sine[24288]=34;
sine[24289]=34;
sine[24290]=34;
sine[24291]=34;
sine[24292]=34;
sine[24293]=34;
sine[24294]=34;
sine[24295]=33;
sine[24296]=33;
sine[24297]=33;
sine[24298]=33;
sine[24299]=33;
sine[24300]=33;
sine[24301]=33;
sine[24302]=33;
sine[24303]=33;
sine[24304]=33;
sine[24305]=33;
sine[24306]=33;
sine[24307]=33;
sine[24308]=33;
sine[24309]=33;
sine[24310]=33;
sine[24311]=33;
sine[24312]=33;
sine[24313]=33;
sine[24314]=33;
sine[24315]=33;
sine[24316]=33;
sine[24317]=33;
sine[24318]=32;
sine[24319]=32;
sine[24320]=32;
sine[24321]=32;
sine[24322]=32;
sine[24323]=32;
sine[24324]=32;
sine[24325]=32;
sine[24326]=32;
sine[24327]=32;
sine[24328]=32;
sine[24329]=32;
sine[24330]=32;
sine[24331]=32;
sine[24332]=32;
sine[24333]=32;
sine[24334]=32;
sine[24335]=32;
sine[24336]=32;
sine[24337]=32;
sine[24338]=32;
sine[24339]=32;
sine[24340]=31;
sine[24341]=31;
sine[24342]=31;
sine[24343]=31;
sine[24344]=31;
sine[24345]=31;
sine[24346]=31;
sine[24347]=31;
sine[24348]=31;
sine[24349]=31;
sine[24350]=31;
sine[24351]=31;
sine[24352]=31;
sine[24353]=31;
sine[24354]=31;
sine[24355]=31;
sine[24356]=31;
sine[24357]=31;
sine[24358]=31;
sine[24359]=31;
sine[24360]=31;
sine[24361]=31;
sine[24362]=30;
sine[24363]=30;
sine[24364]=30;
sine[24365]=30;
sine[24366]=30;
sine[24367]=30;
sine[24368]=30;
sine[24369]=30;
sine[24370]=30;
sine[24371]=30;
sine[24372]=30;
sine[24373]=30;
sine[24374]=30;
sine[24375]=30;
sine[24376]=30;
sine[24377]=30;
sine[24378]=30;
sine[24379]=30;
sine[24380]=30;
sine[24381]=30;
sine[24382]=30;
sine[24383]=30;
sine[24384]=29;
sine[24385]=29;
sine[24386]=29;
sine[24387]=29;
sine[24388]=29;
sine[24389]=29;
sine[24390]=29;
sine[24391]=29;
sine[24392]=29;
sine[24393]=29;
sine[24394]=29;
sine[24395]=29;
sine[24396]=29;
sine[24397]=29;
sine[24398]=29;
sine[24399]=29;
sine[24400]=29;
sine[24401]=29;
sine[24402]=29;
sine[24403]=29;
sine[24404]=29;
sine[24405]=29;
sine[24406]=28;
sine[24407]=28;
sine[24408]=28;
sine[24409]=28;
sine[24410]=28;
sine[24411]=28;
sine[24412]=28;
sine[24413]=28;
sine[24414]=28;
sine[24415]=28;
sine[24416]=28;
sine[24417]=28;
sine[24418]=28;
sine[24419]=28;
sine[24420]=28;
sine[24421]=28;
sine[24422]=28;
sine[24423]=28;
sine[24424]=28;
sine[24425]=28;
sine[24426]=28;
sine[24427]=28;
sine[24428]=27;
sine[24429]=27;
sine[24430]=27;
sine[24431]=27;
sine[24432]=27;
sine[24433]=27;
sine[24434]=27;
sine[24435]=27;
sine[24436]=27;
sine[24437]=27;
sine[24438]=27;
sine[24439]=27;
sine[24440]=27;
sine[24441]=27;
sine[24442]=27;
sine[24443]=27;
sine[24444]=27;
sine[24445]=27;
sine[24446]=27;
sine[24447]=27;
sine[24448]=27;
sine[24449]=27;
sine[24450]=26;
sine[24451]=26;
sine[24452]=26;
sine[24453]=26;
sine[24454]=26;
sine[24455]=26;
sine[24456]=26;
sine[24457]=26;
sine[24458]=26;
sine[24459]=26;
sine[24460]=26;
sine[24461]=26;
sine[24462]=26;
sine[24463]=26;
sine[24464]=26;
sine[24465]=26;
sine[24466]=26;
sine[24467]=26;
sine[24468]=26;
sine[24469]=26;
sine[24470]=26;
sine[24471]=25;
sine[24472]=25;
sine[24473]=25;
sine[24474]=25;
sine[24475]=25;
sine[24476]=25;
sine[24477]=25;
sine[24478]=25;
sine[24479]=25;
sine[24480]=25;
sine[24481]=25;
sine[24482]=25;
sine[24483]=25;
sine[24484]=25;
sine[24485]=25;
sine[24486]=25;
sine[24487]=25;
sine[24488]=25;
sine[24489]=25;
sine[24490]=25;
sine[24491]=25;
sine[24492]=25;
sine[24493]=24;
sine[24494]=24;
sine[24495]=24;
sine[24496]=24;
sine[24497]=24;
sine[24498]=24;
sine[24499]=24;
sine[24500]=24;
sine[24501]=24;
sine[24502]=24;
sine[24503]=24;
sine[24504]=24;
sine[24505]=24;
sine[24506]=24;
sine[24507]=24;
sine[24508]=24;
sine[24509]=24;
sine[24510]=24;
sine[24511]=24;
sine[24512]=24;
sine[24513]=24;
sine[24514]=23;
sine[24515]=23;
sine[24516]=23;
sine[24517]=23;
sine[24518]=23;
sine[24519]=23;
sine[24520]=23;
sine[24521]=23;
sine[24522]=23;
sine[24523]=23;
sine[24524]=23;
sine[24525]=23;
sine[24526]=23;
sine[24527]=23;
sine[24528]=23;
sine[24529]=23;
sine[24530]=23;
sine[24531]=23;
sine[24532]=23;
sine[24533]=23;
sine[24534]=23;
sine[24535]=23;
sine[24536]=22;
sine[24537]=22;
sine[24538]=22;
sine[24539]=22;
sine[24540]=22;
sine[24541]=22;
sine[24542]=22;
sine[24543]=22;
sine[24544]=22;
sine[24545]=22;
sine[24546]=22;
sine[24547]=22;
sine[24548]=22;
sine[24549]=22;
sine[24550]=22;
sine[24551]=22;
sine[24552]=22;
sine[24553]=22;
sine[24554]=22;
sine[24555]=22;
sine[24556]=22;
sine[24557]=21;
sine[24558]=21;
sine[24559]=21;
sine[24560]=21;
sine[24561]=21;
sine[24562]=21;
sine[24563]=21;
sine[24564]=21;
sine[24565]=21;
sine[24566]=21;
sine[24567]=21;
sine[24568]=21;
sine[24569]=21;
sine[24570]=21;
sine[24571]=21;
sine[24572]=21;
sine[24573]=21;
sine[24574]=21;
sine[24575]=21;
sine[24576]=21;
sine[24577]=21;
sine[24578]=20;
sine[24579]=20;
sine[24580]=20;
sine[24581]=20;
sine[24582]=20;
sine[24583]=20;
sine[24584]=20;
sine[24585]=20;
sine[24586]=20;
sine[24587]=20;
sine[24588]=20;
sine[24589]=20;
sine[24590]=20;
sine[24591]=20;
sine[24592]=20;
sine[24593]=20;
sine[24594]=20;
sine[24595]=20;
sine[24596]=20;
sine[24597]=20;
sine[24598]=20;
sine[24599]=19;
sine[24600]=19;
sine[24601]=19;
sine[24602]=19;
sine[24603]=19;
sine[24604]=19;
sine[24605]=19;
sine[24606]=19;
sine[24607]=19;
sine[24608]=19;
sine[24609]=19;
sine[24610]=19;
sine[24611]=19;
sine[24612]=19;
sine[24613]=19;
sine[24614]=19;
sine[24615]=19;
sine[24616]=19;
sine[24617]=19;
sine[24618]=19;
sine[24619]=19;
sine[24620]=18;
sine[24621]=18;
sine[24622]=18;
sine[24623]=18;
sine[24624]=18;
sine[24625]=18;
sine[24626]=18;
sine[24627]=18;
sine[24628]=18;
sine[24629]=18;
sine[24630]=18;
sine[24631]=18;
sine[24632]=18;
sine[24633]=18;
sine[24634]=18;
sine[24635]=18;
sine[24636]=18;
sine[24637]=18;
sine[24638]=18;
sine[24639]=18;
sine[24640]=18;
sine[24641]=17;
sine[24642]=17;
sine[24643]=17;
sine[24644]=17;
sine[24645]=17;
sine[24646]=17;
sine[24647]=17;
sine[24648]=17;
sine[24649]=17;
sine[24650]=17;
sine[24651]=17;
sine[24652]=17;
sine[24653]=17;
sine[24654]=17;
sine[24655]=17;
sine[24656]=17;
sine[24657]=17;
sine[24658]=17;
sine[24659]=17;
sine[24660]=17;
sine[24661]=17;
sine[24662]=16;
sine[24663]=16;
sine[24664]=16;
sine[24665]=16;
sine[24666]=16;
sine[24667]=16;
sine[24668]=16;
sine[24669]=16;
sine[24670]=16;
sine[24671]=16;
sine[24672]=16;
sine[24673]=16;
sine[24674]=16;
sine[24675]=16;
sine[24676]=16;
sine[24677]=16;
sine[24678]=16;
sine[24679]=16;
sine[24680]=16;
sine[24681]=16;
sine[24682]=16;
sine[24683]=15;
sine[24684]=15;
sine[24685]=15;
sine[24686]=15;
sine[24687]=15;
sine[24688]=15;
sine[24689]=15;
sine[24690]=15;
sine[24691]=15;
sine[24692]=15;
sine[24693]=15;
sine[24694]=15;
sine[24695]=15;
sine[24696]=15;
sine[24697]=15;
sine[24698]=15;
sine[24699]=15;
sine[24700]=15;
sine[24701]=15;
sine[24702]=15;
sine[24703]=14;
sine[24704]=14;
sine[24705]=14;
sine[24706]=14;
sine[24707]=14;
sine[24708]=14;
sine[24709]=14;
sine[24710]=14;
sine[24711]=14;
sine[24712]=14;
sine[24713]=14;
sine[24714]=14;
sine[24715]=14;
sine[24716]=14;
sine[24717]=14;
sine[24718]=14;
sine[24719]=14;
sine[24720]=14;
sine[24721]=14;
sine[24722]=14;
sine[24723]=14;
sine[24724]=13;
sine[24725]=13;
sine[24726]=13;
sine[24727]=13;
sine[24728]=13;
sine[24729]=13;
sine[24730]=13;
sine[24731]=13;
sine[24732]=13;
sine[24733]=13;
sine[24734]=13;
sine[24735]=13;
sine[24736]=13;
sine[24737]=13;
sine[24738]=13;
sine[24739]=13;
sine[24740]=13;
sine[24741]=13;
sine[24742]=13;
sine[24743]=13;
sine[24744]=13;
sine[24745]=12;
sine[24746]=12;
sine[24747]=12;
sine[24748]=12;
sine[24749]=12;
sine[24750]=12;
sine[24751]=12;
sine[24752]=12;
sine[24753]=12;
sine[24754]=12;
sine[24755]=12;
sine[24756]=12;
sine[24757]=12;
sine[24758]=12;
sine[24759]=12;
sine[24760]=12;
sine[24761]=12;
sine[24762]=12;
sine[24763]=12;
sine[24764]=12;
sine[24765]=11;
sine[24766]=11;
sine[24767]=11;
sine[24768]=11;
sine[24769]=11;
sine[24770]=11;
sine[24771]=11;
sine[24772]=11;
sine[24773]=11;
sine[24774]=11;
sine[24775]=11;
sine[24776]=11;
sine[24777]=11;
sine[24778]=11;
sine[24779]=11;
sine[24780]=11;
sine[24781]=11;
sine[24782]=11;
sine[24783]=11;
sine[24784]=11;
sine[24785]=11;
sine[24786]=10;
sine[24787]=10;
sine[24788]=10;
sine[24789]=10;
sine[24790]=10;
sine[24791]=10;
sine[24792]=10;
sine[24793]=10;
sine[24794]=10;
sine[24795]=10;
sine[24796]=10;
sine[24797]=10;
sine[24798]=10;
sine[24799]=10;
sine[24800]=10;
sine[24801]=10;
sine[24802]=10;
sine[24803]=10;
sine[24804]=10;
sine[24805]=10;
sine[24806]=9;
sine[24807]=9;
sine[24808]=9;
sine[24809]=9;
sine[24810]=9;
sine[24811]=9;
sine[24812]=9;
sine[24813]=9;
sine[24814]=9;
sine[24815]=9;
sine[24816]=9;
sine[24817]=9;
sine[24818]=9;
sine[24819]=9;
sine[24820]=9;
sine[24821]=9;
sine[24822]=9;
sine[24823]=9;
sine[24824]=9;
sine[24825]=9;
sine[24826]=9;
sine[24827]=8;
sine[24828]=8;
sine[24829]=8;
sine[24830]=8;
sine[24831]=8;
sine[24832]=8;
sine[24833]=8;
sine[24834]=8;
sine[24835]=8;
sine[24836]=8;
sine[24837]=8;
sine[24838]=8;
sine[24839]=8;
sine[24840]=8;
sine[24841]=8;
sine[24842]=8;
sine[24843]=8;
sine[24844]=8;
sine[24845]=8;
sine[24846]=8;
sine[24847]=7;
sine[24848]=7;
sine[24849]=7;
sine[24850]=7;
sine[24851]=7;
sine[24852]=7;
sine[24853]=7;
sine[24854]=7;
sine[24855]=7;
sine[24856]=7;
sine[24857]=7;
sine[24858]=7;
sine[24859]=7;
sine[24860]=7;
sine[24861]=7;
sine[24862]=7;
sine[24863]=7;
sine[24864]=7;
sine[24865]=7;
sine[24866]=7;
sine[24867]=7;
sine[24868]=6;
sine[24869]=6;
sine[24870]=6;
sine[24871]=6;
sine[24872]=6;
sine[24873]=6;
sine[24874]=6;
sine[24875]=6;
sine[24876]=6;
sine[24877]=6;
sine[24878]=6;
sine[24879]=6;
sine[24880]=6;
sine[24881]=6;
sine[24882]=6;
sine[24883]=6;
sine[24884]=6;
sine[24885]=6;
sine[24886]=6;
sine[24887]=6;
sine[24888]=5;
sine[24889]=5;
sine[24890]=5;
sine[24891]=5;
sine[24892]=5;
sine[24893]=5;
sine[24894]=5;
sine[24895]=5;
sine[24896]=5;
sine[24897]=5;
sine[24898]=5;
sine[24899]=5;
sine[24900]=5;
sine[24901]=5;
sine[24902]=5;
sine[24903]=5;
sine[24904]=5;
sine[24905]=5;
sine[24906]=5;
sine[24907]=5;
sine[24908]=5;
sine[24909]=4;
sine[24910]=4;
sine[24911]=4;
sine[24912]=4;
sine[24913]=4;
sine[24914]=4;
sine[24915]=4;
sine[24916]=4;
sine[24917]=4;
sine[24918]=4;
sine[24919]=4;
sine[24920]=4;
sine[24921]=4;
sine[24922]=4;
sine[24923]=4;
sine[24924]=4;
sine[24925]=4;
sine[24926]=4;
sine[24927]=4;
sine[24928]=4;
sine[24929]=3;
sine[24930]=3;
sine[24931]=3;
sine[24932]=3;
sine[24933]=3;
sine[24934]=3;
sine[24935]=3;
sine[24936]=3;
sine[24937]=3;
sine[24938]=3;
sine[24939]=3;
sine[24940]=3;
sine[24941]=3;
sine[24942]=3;
sine[24943]=3;
sine[24944]=3;
sine[24945]=3;
sine[24946]=3;
sine[24947]=3;
sine[24948]=3;
sine[24949]=3;
sine[24950]=2;
sine[24951]=2;
sine[24952]=2;
sine[24953]=2;
sine[24954]=2;
sine[24955]=2;
sine[24956]=2;
sine[24957]=2;
sine[24958]=2;
sine[24959]=2;
sine[24960]=2;
sine[24961]=2;
sine[24962]=2;
sine[24963]=2;
sine[24964]=2;
sine[24965]=2;
sine[24966]=2;
sine[24967]=2;
sine[24968]=2;
sine[24969]=2;
sine[24970]=1;
sine[24971]=1;
sine[24972]=1;
sine[24973]=1;
sine[24974]=1;
sine[24975]=1;
sine[24976]=1;
sine[24977]=1;
sine[24978]=1;
sine[24979]=1;
sine[24980]=1;
sine[24981]=1;
sine[24982]=1;
sine[24983]=1;
sine[24984]=1;
sine[24985]=1;
sine[24986]=1;
sine[24987]=1;
sine[24988]=1;
sine[24989]=1;
sine[24990]=0;
sine[24991]=0;
sine[24992]=0;
sine[24993]=0;
sine[24994]=0;
sine[24995]=0;
sine[24996]=0;
sine[24997]=0;
sine[24998]=0;
sine[24999]=0;
sine[25000]=0;
sine[25001]=0;
sine[25002]=0;
sine[25003]=0;
sine[25004]=0;
sine[25005]=0;
sine[25006]=0;
sine[25007]=0;
sine[25008]=0;
sine[25009]=0;
sine[25010]=0;
sine[25011]=-1;
sine[25012]=-1;
sine[25013]=-1;
sine[25014]=-1;
sine[25015]=-1;
sine[25016]=-1;
sine[25017]=-1;
sine[25018]=-1;
sine[25019]=-1;
sine[25020]=-1;
sine[25021]=-1;
sine[25022]=-1;
sine[25023]=-1;
sine[25024]=-1;
sine[25025]=-1;
sine[25026]=-1;
sine[25027]=-1;
sine[25028]=-1;
sine[25029]=-1;
sine[25030]=-1;
sine[25031]=-2;
sine[25032]=-2;
sine[25033]=-2;
sine[25034]=-2;
sine[25035]=-2;
sine[25036]=-2;
sine[25037]=-2;
sine[25038]=-2;
sine[25039]=-2;
sine[25040]=-2;
sine[25041]=-2;
sine[25042]=-2;
sine[25043]=-2;
sine[25044]=-2;
sine[25045]=-2;
sine[25046]=-2;
sine[25047]=-2;
sine[25048]=-2;
sine[25049]=-2;
sine[25050]=-2;
sine[25051]=-3;
sine[25052]=-3;
sine[25053]=-3;
sine[25054]=-3;
sine[25055]=-3;
sine[25056]=-3;
sine[25057]=-3;
sine[25058]=-3;
sine[25059]=-3;
sine[25060]=-3;
sine[25061]=-3;
sine[25062]=-3;
sine[25063]=-3;
sine[25064]=-3;
sine[25065]=-3;
sine[25066]=-3;
sine[25067]=-3;
sine[25068]=-3;
sine[25069]=-3;
sine[25070]=-3;
sine[25071]=-3;
sine[25072]=-4;
sine[25073]=-4;
sine[25074]=-4;
sine[25075]=-4;
sine[25076]=-4;
sine[25077]=-4;
sine[25078]=-4;
sine[25079]=-4;
sine[25080]=-4;
sine[25081]=-4;
sine[25082]=-4;
sine[25083]=-4;
sine[25084]=-4;
sine[25085]=-4;
sine[25086]=-4;
sine[25087]=-4;
sine[25088]=-4;
sine[25089]=-4;
sine[25090]=-4;
sine[25091]=-4;
sine[25092]=-5;
sine[25093]=-5;
sine[25094]=-5;
sine[25095]=-5;
sine[25096]=-5;
sine[25097]=-5;
sine[25098]=-5;
sine[25099]=-5;
sine[25100]=-5;
sine[25101]=-5;
sine[25102]=-5;
sine[25103]=-5;
sine[25104]=-5;
sine[25105]=-5;
sine[25106]=-5;
sine[25107]=-5;
sine[25108]=-5;
sine[25109]=-5;
sine[25110]=-5;
sine[25111]=-5;
sine[25112]=-5;
sine[25113]=-6;
sine[25114]=-6;
sine[25115]=-6;
sine[25116]=-6;
sine[25117]=-6;
sine[25118]=-6;
sine[25119]=-6;
sine[25120]=-6;
sine[25121]=-6;
sine[25122]=-6;
sine[25123]=-6;
sine[25124]=-6;
sine[25125]=-6;
sine[25126]=-6;
sine[25127]=-6;
sine[25128]=-6;
sine[25129]=-6;
sine[25130]=-6;
sine[25131]=-6;
sine[25132]=-6;
sine[25133]=-7;
sine[25134]=-7;
sine[25135]=-7;
sine[25136]=-7;
sine[25137]=-7;
sine[25138]=-7;
sine[25139]=-7;
sine[25140]=-7;
sine[25141]=-7;
sine[25142]=-7;
sine[25143]=-7;
sine[25144]=-7;
sine[25145]=-7;
sine[25146]=-7;
sine[25147]=-7;
sine[25148]=-7;
sine[25149]=-7;
sine[25150]=-7;
sine[25151]=-7;
sine[25152]=-7;
sine[25153]=-7;
sine[25154]=-8;
sine[25155]=-8;
sine[25156]=-8;
sine[25157]=-8;
sine[25158]=-8;
sine[25159]=-8;
sine[25160]=-8;
sine[25161]=-8;
sine[25162]=-8;
sine[25163]=-8;
sine[25164]=-8;
sine[25165]=-8;
sine[25166]=-8;
sine[25167]=-8;
sine[25168]=-8;
sine[25169]=-8;
sine[25170]=-8;
sine[25171]=-8;
sine[25172]=-8;
sine[25173]=-8;
sine[25174]=-9;
sine[25175]=-9;
sine[25176]=-9;
sine[25177]=-9;
sine[25178]=-9;
sine[25179]=-9;
sine[25180]=-9;
sine[25181]=-9;
sine[25182]=-9;
sine[25183]=-9;
sine[25184]=-9;
sine[25185]=-9;
sine[25186]=-9;
sine[25187]=-9;
sine[25188]=-9;
sine[25189]=-9;
sine[25190]=-9;
sine[25191]=-9;
sine[25192]=-9;
sine[25193]=-9;
sine[25194]=-9;
sine[25195]=-10;
sine[25196]=-10;
sine[25197]=-10;
sine[25198]=-10;
sine[25199]=-10;
sine[25200]=-10;
sine[25201]=-10;
sine[25202]=-10;
sine[25203]=-10;
sine[25204]=-10;
sine[25205]=-10;
sine[25206]=-10;
sine[25207]=-10;
sine[25208]=-10;
sine[25209]=-10;
sine[25210]=-10;
sine[25211]=-10;
sine[25212]=-10;
sine[25213]=-10;
sine[25214]=-10;
sine[25215]=-11;
sine[25216]=-11;
sine[25217]=-11;
sine[25218]=-11;
sine[25219]=-11;
sine[25220]=-11;
sine[25221]=-11;
sine[25222]=-11;
sine[25223]=-11;
sine[25224]=-11;
sine[25225]=-11;
sine[25226]=-11;
sine[25227]=-11;
sine[25228]=-11;
sine[25229]=-11;
sine[25230]=-11;
sine[25231]=-11;
sine[25232]=-11;
sine[25233]=-11;
sine[25234]=-11;
sine[25235]=-11;
sine[25236]=-12;
sine[25237]=-12;
sine[25238]=-12;
sine[25239]=-12;
sine[25240]=-12;
sine[25241]=-12;
sine[25242]=-12;
sine[25243]=-12;
sine[25244]=-12;
sine[25245]=-12;
sine[25246]=-12;
sine[25247]=-12;
sine[25248]=-12;
sine[25249]=-12;
sine[25250]=-12;
sine[25251]=-12;
sine[25252]=-12;
sine[25253]=-12;
sine[25254]=-12;
sine[25255]=-12;
sine[25256]=-13;
sine[25257]=-13;
sine[25258]=-13;
sine[25259]=-13;
sine[25260]=-13;
sine[25261]=-13;
sine[25262]=-13;
sine[25263]=-13;
sine[25264]=-13;
sine[25265]=-13;
sine[25266]=-13;
sine[25267]=-13;
sine[25268]=-13;
sine[25269]=-13;
sine[25270]=-13;
sine[25271]=-13;
sine[25272]=-13;
sine[25273]=-13;
sine[25274]=-13;
sine[25275]=-13;
sine[25276]=-13;
sine[25277]=-14;
sine[25278]=-14;
sine[25279]=-14;
sine[25280]=-14;
sine[25281]=-14;
sine[25282]=-14;
sine[25283]=-14;
sine[25284]=-14;
sine[25285]=-14;
sine[25286]=-14;
sine[25287]=-14;
sine[25288]=-14;
sine[25289]=-14;
sine[25290]=-14;
sine[25291]=-14;
sine[25292]=-14;
sine[25293]=-14;
sine[25294]=-14;
sine[25295]=-14;
sine[25296]=-14;
sine[25297]=-14;
sine[25298]=-15;
sine[25299]=-15;
sine[25300]=-15;
sine[25301]=-15;
sine[25302]=-15;
sine[25303]=-15;
sine[25304]=-15;
sine[25305]=-15;
sine[25306]=-15;
sine[25307]=-15;
sine[25308]=-15;
sine[25309]=-15;
sine[25310]=-15;
sine[25311]=-15;
sine[25312]=-15;
sine[25313]=-15;
sine[25314]=-15;
sine[25315]=-15;
sine[25316]=-15;
sine[25317]=-15;
sine[25318]=-16;
sine[25319]=-16;
sine[25320]=-16;
sine[25321]=-16;
sine[25322]=-16;
sine[25323]=-16;
sine[25324]=-16;
sine[25325]=-16;
sine[25326]=-16;
sine[25327]=-16;
sine[25328]=-16;
sine[25329]=-16;
sine[25330]=-16;
sine[25331]=-16;
sine[25332]=-16;
sine[25333]=-16;
sine[25334]=-16;
sine[25335]=-16;
sine[25336]=-16;
sine[25337]=-16;
sine[25338]=-16;
sine[25339]=-17;
sine[25340]=-17;
sine[25341]=-17;
sine[25342]=-17;
sine[25343]=-17;
sine[25344]=-17;
sine[25345]=-17;
sine[25346]=-17;
sine[25347]=-17;
sine[25348]=-17;
sine[25349]=-17;
sine[25350]=-17;
sine[25351]=-17;
sine[25352]=-17;
sine[25353]=-17;
sine[25354]=-17;
sine[25355]=-17;
sine[25356]=-17;
sine[25357]=-17;
sine[25358]=-17;
sine[25359]=-17;
sine[25360]=-18;
sine[25361]=-18;
sine[25362]=-18;
sine[25363]=-18;
sine[25364]=-18;
sine[25365]=-18;
sine[25366]=-18;
sine[25367]=-18;
sine[25368]=-18;
sine[25369]=-18;
sine[25370]=-18;
sine[25371]=-18;
sine[25372]=-18;
sine[25373]=-18;
sine[25374]=-18;
sine[25375]=-18;
sine[25376]=-18;
sine[25377]=-18;
sine[25378]=-18;
sine[25379]=-18;
sine[25380]=-18;
sine[25381]=-19;
sine[25382]=-19;
sine[25383]=-19;
sine[25384]=-19;
sine[25385]=-19;
sine[25386]=-19;
sine[25387]=-19;
sine[25388]=-19;
sine[25389]=-19;
sine[25390]=-19;
sine[25391]=-19;
sine[25392]=-19;
sine[25393]=-19;
sine[25394]=-19;
sine[25395]=-19;
sine[25396]=-19;
sine[25397]=-19;
sine[25398]=-19;
sine[25399]=-19;
sine[25400]=-19;
sine[25401]=-19;
sine[25402]=-20;
sine[25403]=-20;
sine[25404]=-20;
sine[25405]=-20;
sine[25406]=-20;
sine[25407]=-20;
sine[25408]=-20;
sine[25409]=-20;
sine[25410]=-20;
sine[25411]=-20;
sine[25412]=-20;
sine[25413]=-20;
sine[25414]=-20;
sine[25415]=-20;
sine[25416]=-20;
sine[25417]=-20;
sine[25418]=-20;
sine[25419]=-20;
sine[25420]=-20;
sine[25421]=-20;
sine[25422]=-20;
sine[25423]=-21;
sine[25424]=-21;
sine[25425]=-21;
sine[25426]=-21;
sine[25427]=-21;
sine[25428]=-21;
sine[25429]=-21;
sine[25430]=-21;
sine[25431]=-21;
sine[25432]=-21;
sine[25433]=-21;
sine[25434]=-21;
sine[25435]=-21;
sine[25436]=-21;
sine[25437]=-21;
sine[25438]=-21;
sine[25439]=-21;
sine[25440]=-21;
sine[25441]=-21;
sine[25442]=-21;
sine[25443]=-21;
sine[25444]=-22;
sine[25445]=-22;
sine[25446]=-22;
sine[25447]=-22;
sine[25448]=-22;
sine[25449]=-22;
sine[25450]=-22;
sine[25451]=-22;
sine[25452]=-22;
sine[25453]=-22;
sine[25454]=-22;
sine[25455]=-22;
sine[25456]=-22;
sine[25457]=-22;
sine[25458]=-22;
sine[25459]=-22;
sine[25460]=-22;
sine[25461]=-22;
sine[25462]=-22;
sine[25463]=-22;
sine[25464]=-22;
sine[25465]=-23;
sine[25466]=-23;
sine[25467]=-23;
sine[25468]=-23;
sine[25469]=-23;
sine[25470]=-23;
sine[25471]=-23;
sine[25472]=-23;
sine[25473]=-23;
sine[25474]=-23;
sine[25475]=-23;
sine[25476]=-23;
sine[25477]=-23;
sine[25478]=-23;
sine[25479]=-23;
sine[25480]=-23;
sine[25481]=-23;
sine[25482]=-23;
sine[25483]=-23;
sine[25484]=-23;
sine[25485]=-23;
sine[25486]=-23;
sine[25487]=-24;
sine[25488]=-24;
sine[25489]=-24;
sine[25490]=-24;
sine[25491]=-24;
sine[25492]=-24;
sine[25493]=-24;
sine[25494]=-24;
sine[25495]=-24;
sine[25496]=-24;
sine[25497]=-24;
sine[25498]=-24;
sine[25499]=-24;
sine[25500]=-24;
sine[25501]=-24;
sine[25502]=-24;
sine[25503]=-24;
sine[25504]=-24;
sine[25505]=-24;
sine[25506]=-24;
sine[25507]=-24;
sine[25508]=-25;
sine[25509]=-25;
sine[25510]=-25;
sine[25511]=-25;
sine[25512]=-25;
sine[25513]=-25;
sine[25514]=-25;
sine[25515]=-25;
sine[25516]=-25;
sine[25517]=-25;
sine[25518]=-25;
sine[25519]=-25;
sine[25520]=-25;
sine[25521]=-25;
sine[25522]=-25;
sine[25523]=-25;
sine[25524]=-25;
sine[25525]=-25;
sine[25526]=-25;
sine[25527]=-25;
sine[25528]=-25;
sine[25529]=-25;
sine[25530]=-26;
sine[25531]=-26;
sine[25532]=-26;
sine[25533]=-26;
sine[25534]=-26;
sine[25535]=-26;
sine[25536]=-26;
sine[25537]=-26;
sine[25538]=-26;
sine[25539]=-26;
sine[25540]=-26;
sine[25541]=-26;
sine[25542]=-26;
sine[25543]=-26;
sine[25544]=-26;
sine[25545]=-26;
sine[25546]=-26;
sine[25547]=-26;
sine[25548]=-26;
sine[25549]=-26;
sine[25550]=-26;
sine[25551]=-27;
sine[25552]=-27;
sine[25553]=-27;
sine[25554]=-27;
sine[25555]=-27;
sine[25556]=-27;
sine[25557]=-27;
sine[25558]=-27;
sine[25559]=-27;
sine[25560]=-27;
sine[25561]=-27;
sine[25562]=-27;
sine[25563]=-27;
sine[25564]=-27;
sine[25565]=-27;
sine[25566]=-27;
sine[25567]=-27;
sine[25568]=-27;
sine[25569]=-27;
sine[25570]=-27;
sine[25571]=-27;
sine[25572]=-27;
sine[25573]=-28;
sine[25574]=-28;
sine[25575]=-28;
sine[25576]=-28;
sine[25577]=-28;
sine[25578]=-28;
sine[25579]=-28;
sine[25580]=-28;
sine[25581]=-28;
sine[25582]=-28;
sine[25583]=-28;
sine[25584]=-28;
sine[25585]=-28;
sine[25586]=-28;
sine[25587]=-28;
sine[25588]=-28;
sine[25589]=-28;
sine[25590]=-28;
sine[25591]=-28;
sine[25592]=-28;
sine[25593]=-28;
sine[25594]=-28;
sine[25595]=-29;
sine[25596]=-29;
sine[25597]=-29;
sine[25598]=-29;
sine[25599]=-29;
sine[25600]=-29;
sine[25601]=-29;
sine[25602]=-29;
sine[25603]=-29;
sine[25604]=-29;
sine[25605]=-29;
sine[25606]=-29;
sine[25607]=-29;
sine[25608]=-29;
sine[25609]=-29;
sine[25610]=-29;
sine[25611]=-29;
sine[25612]=-29;
sine[25613]=-29;
sine[25614]=-29;
sine[25615]=-29;
sine[25616]=-29;
sine[25617]=-30;
sine[25618]=-30;
sine[25619]=-30;
sine[25620]=-30;
sine[25621]=-30;
sine[25622]=-30;
sine[25623]=-30;
sine[25624]=-30;
sine[25625]=-30;
sine[25626]=-30;
sine[25627]=-30;
sine[25628]=-30;
sine[25629]=-30;
sine[25630]=-30;
sine[25631]=-30;
sine[25632]=-30;
sine[25633]=-30;
sine[25634]=-30;
sine[25635]=-30;
sine[25636]=-30;
sine[25637]=-30;
sine[25638]=-30;
sine[25639]=-31;
sine[25640]=-31;
sine[25641]=-31;
sine[25642]=-31;
sine[25643]=-31;
sine[25644]=-31;
sine[25645]=-31;
sine[25646]=-31;
sine[25647]=-31;
sine[25648]=-31;
sine[25649]=-31;
sine[25650]=-31;
sine[25651]=-31;
sine[25652]=-31;
sine[25653]=-31;
sine[25654]=-31;
sine[25655]=-31;
sine[25656]=-31;
sine[25657]=-31;
sine[25658]=-31;
sine[25659]=-31;
sine[25660]=-31;
sine[25661]=-32;
sine[25662]=-32;
sine[25663]=-32;
sine[25664]=-32;
sine[25665]=-32;
sine[25666]=-32;
sine[25667]=-32;
sine[25668]=-32;
sine[25669]=-32;
sine[25670]=-32;
sine[25671]=-32;
sine[25672]=-32;
sine[25673]=-32;
sine[25674]=-32;
sine[25675]=-32;
sine[25676]=-32;
sine[25677]=-32;
sine[25678]=-32;
sine[25679]=-32;
sine[25680]=-32;
sine[25681]=-32;
sine[25682]=-32;
sine[25683]=-33;
sine[25684]=-33;
sine[25685]=-33;
sine[25686]=-33;
sine[25687]=-33;
sine[25688]=-33;
sine[25689]=-33;
sine[25690]=-33;
sine[25691]=-33;
sine[25692]=-33;
sine[25693]=-33;
sine[25694]=-33;
sine[25695]=-33;
sine[25696]=-33;
sine[25697]=-33;
sine[25698]=-33;
sine[25699]=-33;
sine[25700]=-33;
sine[25701]=-33;
sine[25702]=-33;
sine[25703]=-33;
sine[25704]=-33;
sine[25705]=-33;
sine[25706]=-34;
sine[25707]=-34;
sine[25708]=-34;
sine[25709]=-34;
sine[25710]=-34;
sine[25711]=-34;
sine[25712]=-34;
sine[25713]=-34;
sine[25714]=-34;
sine[25715]=-34;
sine[25716]=-34;
sine[25717]=-34;
sine[25718]=-34;
sine[25719]=-34;
sine[25720]=-34;
sine[25721]=-34;
sine[25722]=-34;
sine[25723]=-34;
sine[25724]=-34;
sine[25725]=-34;
sine[25726]=-34;
sine[25727]=-34;
sine[25728]=-35;
sine[25729]=-35;
sine[25730]=-35;
sine[25731]=-35;
sine[25732]=-35;
sine[25733]=-35;
sine[25734]=-35;
sine[25735]=-35;
sine[25736]=-35;
sine[25737]=-35;
sine[25738]=-35;
sine[25739]=-35;
sine[25740]=-35;
sine[25741]=-35;
sine[25742]=-35;
sine[25743]=-35;
sine[25744]=-35;
sine[25745]=-35;
sine[25746]=-35;
sine[25747]=-35;
sine[25748]=-35;
sine[25749]=-35;
sine[25750]=-35;
sine[25751]=-36;
sine[25752]=-36;
sine[25753]=-36;
sine[25754]=-36;
sine[25755]=-36;
sine[25756]=-36;
sine[25757]=-36;
sine[25758]=-36;
sine[25759]=-36;
sine[25760]=-36;
sine[25761]=-36;
sine[25762]=-36;
sine[25763]=-36;
sine[25764]=-36;
sine[25765]=-36;
sine[25766]=-36;
sine[25767]=-36;
sine[25768]=-36;
sine[25769]=-36;
sine[25770]=-36;
sine[25771]=-36;
sine[25772]=-36;
sine[25773]=-36;
sine[25774]=-37;
sine[25775]=-37;
sine[25776]=-37;
sine[25777]=-37;
sine[25778]=-37;
sine[25779]=-37;
sine[25780]=-37;
sine[25781]=-37;
sine[25782]=-37;
sine[25783]=-37;
sine[25784]=-37;
sine[25785]=-37;
sine[25786]=-37;
sine[25787]=-37;
sine[25788]=-37;
sine[25789]=-37;
sine[25790]=-37;
sine[25791]=-37;
sine[25792]=-37;
sine[25793]=-37;
sine[25794]=-37;
sine[25795]=-37;
sine[25796]=-37;
sine[25797]=-38;
sine[25798]=-38;
sine[25799]=-38;
sine[25800]=-38;
sine[25801]=-38;
sine[25802]=-38;
sine[25803]=-38;
sine[25804]=-38;
sine[25805]=-38;
sine[25806]=-38;
sine[25807]=-38;
sine[25808]=-38;
sine[25809]=-38;
sine[25810]=-38;
sine[25811]=-38;
sine[25812]=-38;
sine[25813]=-38;
sine[25814]=-38;
sine[25815]=-38;
sine[25816]=-38;
sine[25817]=-38;
sine[25818]=-38;
sine[25819]=-38;
sine[25820]=-38;
sine[25821]=-39;
sine[25822]=-39;
sine[25823]=-39;
sine[25824]=-39;
sine[25825]=-39;
sine[25826]=-39;
sine[25827]=-39;
sine[25828]=-39;
sine[25829]=-39;
sine[25830]=-39;
sine[25831]=-39;
sine[25832]=-39;
sine[25833]=-39;
sine[25834]=-39;
sine[25835]=-39;
sine[25836]=-39;
sine[25837]=-39;
sine[25838]=-39;
sine[25839]=-39;
sine[25840]=-39;
sine[25841]=-39;
sine[25842]=-39;
sine[25843]=-39;
sine[25844]=-40;
sine[25845]=-40;
sine[25846]=-40;
sine[25847]=-40;
sine[25848]=-40;
sine[25849]=-40;
sine[25850]=-40;
sine[25851]=-40;
sine[25852]=-40;
sine[25853]=-40;
sine[25854]=-40;
sine[25855]=-40;
sine[25856]=-40;
sine[25857]=-40;
sine[25858]=-40;
sine[25859]=-40;
sine[25860]=-40;
sine[25861]=-40;
sine[25862]=-40;
sine[25863]=-40;
sine[25864]=-40;
sine[25865]=-40;
sine[25866]=-40;
sine[25867]=-40;
sine[25868]=-41;
sine[25869]=-41;
sine[25870]=-41;
sine[25871]=-41;
sine[25872]=-41;
sine[25873]=-41;
sine[25874]=-41;
sine[25875]=-41;
sine[25876]=-41;
sine[25877]=-41;
sine[25878]=-41;
sine[25879]=-41;
sine[25880]=-41;
sine[25881]=-41;
sine[25882]=-41;
sine[25883]=-41;
sine[25884]=-41;
sine[25885]=-41;
sine[25886]=-41;
sine[25887]=-41;
sine[25888]=-41;
sine[25889]=-41;
sine[25890]=-41;
sine[25891]=-41;
sine[25892]=-42;
sine[25893]=-42;
sine[25894]=-42;
sine[25895]=-42;
sine[25896]=-42;
sine[25897]=-42;
sine[25898]=-42;
sine[25899]=-42;
sine[25900]=-42;
sine[25901]=-42;
sine[25902]=-42;
sine[25903]=-42;
sine[25904]=-42;
sine[25905]=-42;
sine[25906]=-42;
sine[25907]=-42;
sine[25908]=-42;
sine[25909]=-42;
sine[25910]=-42;
sine[25911]=-42;
sine[25912]=-42;
sine[25913]=-42;
sine[25914]=-42;
sine[25915]=-42;
sine[25916]=-43;
sine[25917]=-43;
sine[25918]=-43;
sine[25919]=-43;
sine[25920]=-43;
sine[25921]=-43;
sine[25922]=-43;
sine[25923]=-43;
sine[25924]=-43;
sine[25925]=-43;
sine[25926]=-43;
sine[25927]=-43;
sine[25928]=-43;
sine[25929]=-43;
sine[25930]=-43;
sine[25931]=-43;
sine[25932]=-43;
sine[25933]=-43;
sine[25934]=-43;
sine[25935]=-43;
sine[25936]=-43;
sine[25937]=-43;
sine[25938]=-43;
sine[25939]=-43;
sine[25940]=-44;
sine[25941]=-44;
sine[25942]=-44;
sine[25943]=-44;
sine[25944]=-44;
sine[25945]=-44;
sine[25946]=-44;
sine[25947]=-44;
sine[25948]=-44;
sine[25949]=-44;
sine[25950]=-44;
sine[25951]=-44;
sine[25952]=-44;
sine[25953]=-44;
sine[25954]=-44;
sine[25955]=-44;
sine[25956]=-44;
sine[25957]=-44;
sine[25958]=-44;
sine[25959]=-44;
sine[25960]=-44;
sine[25961]=-44;
sine[25962]=-44;
sine[25963]=-44;
sine[25964]=-44;
sine[25965]=-45;
sine[25966]=-45;
sine[25967]=-45;
sine[25968]=-45;
sine[25969]=-45;
sine[25970]=-45;
sine[25971]=-45;
sine[25972]=-45;
sine[25973]=-45;
sine[25974]=-45;
sine[25975]=-45;
sine[25976]=-45;
sine[25977]=-45;
sine[25978]=-45;
sine[25979]=-45;
sine[25980]=-45;
sine[25981]=-45;
sine[25982]=-45;
sine[25983]=-45;
sine[25984]=-45;
sine[25985]=-45;
sine[25986]=-45;
sine[25987]=-45;
sine[25988]=-45;
sine[25989]=-45;
sine[25990]=-46;
sine[25991]=-46;
sine[25992]=-46;
sine[25993]=-46;
sine[25994]=-46;
sine[25995]=-46;
sine[25996]=-46;
sine[25997]=-46;
sine[25998]=-46;
sine[25999]=-46;
sine[26000]=-46;
sine[26001]=-46;
sine[26002]=-46;
sine[26003]=-46;
sine[26004]=-46;
sine[26005]=-46;
sine[26006]=-46;
sine[26007]=-46;
sine[26008]=-46;
sine[26009]=-46;
sine[26010]=-46;
sine[26011]=-46;
sine[26012]=-46;
sine[26013]=-46;
sine[26014]=-46;
sine[26015]=-47;
sine[26016]=-47;
sine[26017]=-47;
sine[26018]=-47;
sine[26019]=-47;
sine[26020]=-47;
sine[26021]=-47;
sine[26022]=-47;
sine[26023]=-47;
sine[26024]=-47;
sine[26025]=-47;
sine[26026]=-47;
sine[26027]=-47;
sine[26028]=-47;
sine[26029]=-47;
sine[26030]=-47;
sine[26031]=-47;
sine[26032]=-47;
sine[26033]=-47;
sine[26034]=-47;
sine[26035]=-47;
sine[26036]=-47;
sine[26037]=-47;
sine[26038]=-47;
sine[26039]=-47;
sine[26040]=-47;
sine[26041]=-48;
sine[26042]=-48;
sine[26043]=-48;
sine[26044]=-48;
sine[26045]=-48;
sine[26046]=-48;
sine[26047]=-48;
sine[26048]=-48;
sine[26049]=-48;
sine[26050]=-48;
sine[26051]=-48;
sine[26052]=-48;
sine[26053]=-48;
sine[26054]=-48;
sine[26055]=-48;
sine[26056]=-48;
sine[26057]=-48;
sine[26058]=-48;
sine[26059]=-48;
sine[26060]=-48;
sine[26061]=-48;
sine[26062]=-48;
sine[26063]=-48;
sine[26064]=-48;
sine[26065]=-48;
sine[26066]=-49;
sine[26067]=-49;
sine[26068]=-49;
sine[26069]=-49;
sine[26070]=-49;
sine[26071]=-49;
sine[26072]=-49;
sine[26073]=-49;
sine[26074]=-49;
sine[26075]=-49;
sine[26076]=-49;
sine[26077]=-49;
sine[26078]=-49;
sine[26079]=-49;
sine[26080]=-49;
sine[26081]=-49;
sine[26082]=-49;
sine[26083]=-49;
sine[26084]=-49;
sine[26085]=-49;
sine[26086]=-49;
sine[26087]=-49;
sine[26088]=-49;
sine[26089]=-49;
sine[26090]=-49;
sine[26091]=-49;
sine[26092]=-49;
sine[26093]=-50;
sine[26094]=-50;
sine[26095]=-50;
sine[26096]=-50;
sine[26097]=-50;
sine[26098]=-50;
sine[26099]=-50;
sine[26100]=-50;
sine[26101]=-50;
sine[26102]=-50;
sine[26103]=-50;
sine[26104]=-50;
sine[26105]=-50;
sine[26106]=-50;
sine[26107]=-50;
sine[26108]=-50;
sine[26109]=-50;
sine[26110]=-50;
sine[26111]=-50;
sine[26112]=-50;
sine[26113]=-50;
sine[26114]=-50;
sine[26115]=-50;
sine[26116]=-50;
sine[26117]=-50;
sine[26118]=-50;
sine[26119]=-51;
sine[26120]=-51;
sine[26121]=-51;
sine[26122]=-51;
sine[26123]=-51;
sine[26124]=-51;
sine[26125]=-51;
sine[26126]=-51;
sine[26127]=-51;
sine[26128]=-51;
sine[26129]=-51;
sine[26130]=-51;
sine[26131]=-51;
sine[26132]=-51;
sine[26133]=-51;
sine[26134]=-51;
sine[26135]=-51;
sine[26136]=-51;
sine[26137]=-51;
sine[26138]=-51;
sine[26139]=-51;
sine[26140]=-51;
sine[26141]=-51;
sine[26142]=-51;
sine[26143]=-51;
sine[26144]=-51;
sine[26145]=-51;
sine[26146]=-52;
sine[26147]=-52;
sine[26148]=-52;
sine[26149]=-52;
sine[26150]=-52;
sine[26151]=-52;
sine[26152]=-52;
sine[26153]=-52;
sine[26154]=-52;
sine[26155]=-52;
sine[26156]=-52;
sine[26157]=-52;
sine[26158]=-52;
sine[26159]=-52;
sine[26160]=-52;
sine[26161]=-52;
sine[26162]=-52;
sine[26163]=-52;
sine[26164]=-52;
sine[26165]=-52;
sine[26166]=-52;
sine[26167]=-52;
sine[26168]=-52;
sine[26169]=-52;
sine[26170]=-52;
sine[26171]=-52;
sine[26172]=-52;
sine[26173]=-53;
sine[26174]=-53;
sine[26175]=-53;
sine[26176]=-53;
sine[26177]=-53;
sine[26178]=-53;
sine[26179]=-53;
sine[26180]=-53;
sine[26181]=-53;
sine[26182]=-53;
sine[26183]=-53;
sine[26184]=-53;
sine[26185]=-53;
sine[26186]=-53;
sine[26187]=-53;
sine[26188]=-53;
sine[26189]=-53;
sine[26190]=-53;
sine[26191]=-53;
sine[26192]=-53;
sine[26193]=-53;
sine[26194]=-53;
sine[26195]=-53;
sine[26196]=-53;
sine[26197]=-53;
sine[26198]=-53;
sine[26199]=-53;
sine[26200]=-53;
sine[26201]=-54;
sine[26202]=-54;
sine[26203]=-54;
sine[26204]=-54;
sine[26205]=-54;
sine[26206]=-54;
sine[26207]=-54;
sine[26208]=-54;
sine[26209]=-54;
sine[26210]=-54;
sine[26211]=-54;
sine[26212]=-54;
sine[26213]=-54;
sine[26214]=-54;
sine[26215]=-54;
sine[26216]=-54;
sine[26217]=-54;
sine[26218]=-54;
sine[26219]=-54;
sine[26220]=-54;
sine[26221]=-54;
sine[26222]=-54;
sine[26223]=-54;
sine[26224]=-54;
sine[26225]=-54;
sine[26226]=-54;
sine[26227]=-54;
sine[26228]=-54;
sine[26229]=-55;
sine[26230]=-55;
sine[26231]=-55;
sine[26232]=-55;
sine[26233]=-55;
sine[26234]=-55;
sine[26235]=-55;
sine[26236]=-55;
sine[26237]=-55;
sine[26238]=-55;
sine[26239]=-55;
sine[26240]=-55;
sine[26241]=-55;
sine[26242]=-55;
sine[26243]=-55;
sine[26244]=-55;
sine[26245]=-55;
sine[26246]=-55;
sine[26247]=-55;
sine[26248]=-55;
sine[26249]=-55;
sine[26250]=-55;
sine[26251]=-55;
sine[26252]=-55;
sine[26253]=-55;
sine[26254]=-55;
sine[26255]=-55;
sine[26256]=-55;
sine[26257]=-55;
sine[26258]=-56;
sine[26259]=-56;
sine[26260]=-56;
sine[26261]=-56;
sine[26262]=-56;
sine[26263]=-56;
sine[26264]=-56;
sine[26265]=-56;
sine[26266]=-56;
sine[26267]=-56;
sine[26268]=-56;
sine[26269]=-56;
sine[26270]=-56;
sine[26271]=-56;
sine[26272]=-56;
sine[26273]=-56;
sine[26274]=-56;
sine[26275]=-56;
sine[26276]=-56;
sine[26277]=-56;
sine[26278]=-56;
sine[26279]=-56;
sine[26280]=-56;
sine[26281]=-56;
sine[26282]=-56;
sine[26283]=-56;
sine[26284]=-56;
sine[26285]=-56;
sine[26286]=-56;
sine[26287]=-57;
sine[26288]=-57;
sine[26289]=-57;
sine[26290]=-57;
sine[26291]=-57;
sine[26292]=-57;
sine[26293]=-57;
sine[26294]=-57;
sine[26295]=-57;
sine[26296]=-57;
sine[26297]=-57;
sine[26298]=-57;
sine[26299]=-57;
sine[26300]=-57;
sine[26301]=-57;
sine[26302]=-57;
sine[26303]=-57;
sine[26304]=-57;
sine[26305]=-57;
sine[26306]=-57;
sine[26307]=-57;
sine[26308]=-57;
sine[26309]=-57;
sine[26310]=-57;
sine[26311]=-57;
sine[26312]=-57;
sine[26313]=-57;
sine[26314]=-57;
sine[26315]=-57;
sine[26316]=-57;
sine[26317]=-58;
sine[26318]=-58;
sine[26319]=-58;
sine[26320]=-58;
sine[26321]=-58;
sine[26322]=-58;
sine[26323]=-58;
sine[26324]=-58;
sine[26325]=-58;
sine[26326]=-58;
sine[26327]=-58;
sine[26328]=-58;
sine[26329]=-58;
sine[26330]=-58;
sine[26331]=-58;
sine[26332]=-58;
sine[26333]=-58;
sine[26334]=-58;
sine[26335]=-58;
sine[26336]=-58;
sine[26337]=-58;
sine[26338]=-58;
sine[26339]=-58;
sine[26340]=-58;
sine[26341]=-58;
sine[26342]=-58;
sine[26343]=-58;
sine[26344]=-58;
sine[26345]=-58;
sine[26346]=-58;
sine[26347]=-59;
sine[26348]=-59;
sine[26349]=-59;
sine[26350]=-59;
sine[26351]=-59;
sine[26352]=-59;
sine[26353]=-59;
sine[26354]=-59;
sine[26355]=-59;
sine[26356]=-59;
sine[26357]=-59;
sine[26358]=-59;
sine[26359]=-59;
sine[26360]=-59;
sine[26361]=-59;
sine[26362]=-59;
sine[26363]=-59;
sine[26364]=-59;
sine[26365]=-59;
sine[26366]=-59;
sine[26367]=-59;
sine[26368]=-59;
sine[26369]=-59;
sine[26370]=-59;
sine[26371]=-59;
sine[26372]=-59;
sine[26373]=-59;
sine[26374]=-59;
sine[26375]=-59;
sine[26376]=-59;
sine[26377]=-59;
sine[26378]=-60;
sine[26379]=-60;
sine[26380]=-60;
sine[26381]=-60;
sine[26382]=-60;
sine[26383]=-60;
sine[26384]=-60;
sine[26385]=-60;
sine[26386]=-60;
sine[26387]=-60;
sine[26388]=-60;
sine[26389]=-60;
sine[26390]=-60;
sine[26391]=-60;
sine[26392]=-60;
sine[26393]=-60;
sine[26394]=-60;
sine[26395]=-60;
sine[26396]=-60;
sine[26397]=-60;
sine[26398]=-60;
sine[26399]=-60;
sine[26400]=-60;
sine[26401]=-60;
sine[26402]=-60;
sine[26403]=-60;
sine[26404]=-60;
sine[26405]=-60;
sine[26406]=-60;
sine[26407]=-60;
sine[26408]=-60;
sine[26409]=-60;
sine[26410]=-61;
sine[26411]=-61;
sine[26412]=-61;
sine[26413]=-61;
sine[26414]=-61;
sine[26415]=-61;
sine[26416]=-61;
sine[26417]=-61;
sine[26418]=-61;
sine[26419]=-61;
sine[26420]=-61;
sine[26421]=-61;
sine[26422]=-61;
sine[26423]=-61;
sine[26424]=-61;
sine[26425]=-61;
sine[26426]=-61;
sine[26427]=-61;
sine[26428]=-61;
sine[26429]=-61;
sine[26430]=-61;
sine[26431]=-61;
sine[26432]=-61;
sine[26433]=-61;
sine[26434]=-61;
sine[26435]=-61;
sine[26436]=-61;
sine[26437]=-61;
sine[26438]=-61;
sine[26439]=-61;
sine[26440]=-61;
sine[26441]=-61;
sine[26442]=-61;
sine[26443]=-62;
sine[26444]=-62;
sine[26445]=-62;
sine[26446]=-62;
sine[26447]=-62;
sine[26448]=-62;
sine[26449]=-62;
sine[26450]=-62;
sine[26451]=-62;
sine[26452]=-62;
sine[26453]=-62;
sine[26454]=-62;
sine[26455]=-62;
sine[26456]=-62;
sine[26457]=-62;
sine[26458]=-62;
sine[26459]=-62;
sine[26460]=-62;
sine[26461]=-62;
sine[26462]=-62;
sine[26463]=-62;
sine[26464]=-62;
sine[26465]=-62;
sine[26466]=-62;
sine[26467]=-62;
sine[26468]=-62;
sine[26469]=-62;
sine[26470]=-62;
sine[26471]=-62;
sine[26472]=-62;
sine[26473]=-62;
sine[26474]=-62;
sine[26475]=-62;
sine[26476]=-63;
sine[26477]=-63;
sine[26478]=-63;
sine[26479]=-63;
sine[26480]=-63;
sine[26481]=-63;
sine[26482]=-63;
sine[26483]=-63;
sine[26484]=-63;
sine[26485]=-63;
sine[26486]=-63;
sine[26487]=-63;
sine[26488]=-63;
sine[26489]=-63;
sine[26490]=-63;
sine[26491]=-63;
sine[26492]=-63;
sine[26493]=-63;
sine[26494]=-63;
sine[26495]=-63;
sine[26496]=-63;
sine[26497]=-63;
sine[26498]=-63;
sine[26499]=-63;
sine[26500]=-63;
sine[26501]=-63;
sine[26502]=-63;
sine[26503]=-63;
sine[26504]=-63;
sine[26505]=-63;
sine[26506]=-63;
sine[26507]=-63;
sine[26508]=-63;
sine[26509]=-63;
sine[26510]=-63;
sine[26511]=-64;
sine[26512]=-64;
sine[26513]=-64;
sine[26514]=-64;
sine[26515]=-64;
sine[26516]=-64;
sine[26517]=-64;
sine[26518]=-64;
sine[26519]=-64;
sine[26520]=-64;
sine[26521]=-64;
sine[26522]=-64;
sine[26523]=-64;
sine[26524]=-64;
sine[26525]=-64;
sine[26526]=-64;
sine[26527]=-64;
sine[26528]=-64;
sine[26529]=-64;
sine[26530]=-64;
sine[26531]=-64;
sine[26532]=-64;
sine[26533]=-64;
sine[26534]=-64;
sine[26535]=-64;
sine[26536]=-64;
sine[26537]=-64;
sine[26538]=-64;
sine[26539]=-64;
sine[26540]=-64;
sine[26541]=-64;
sine[26542]=-64;
sine[26543]=-64;
sine[26544]=-64;
sine[26545]=-64;
sine[26546]=-65;
sine[26547]=-65;
sine[26548]=-65;
sine[26549]=-65;
sine[26550]=-65;
sine[26551]=-65;
sine[26552]=-65;
sine[26553]=-65;
sine[26554]=-65;
sine[26555]=-65;
sine[26556]=-65;
sine[26557]=-65;
sine[26558]=-65;
sine[26559]=-65;
sine[26560]=-65;
sine[26561]=-65;
sine[26562]=-65;
sine[26563]=-65;
sine[26564]=-65;
sine[26565]=-65;
sine[26566]=-65;
sine[26567]=-65;
sine[26568]=-65;
sine[26569]=-65;
sine[26570]=-65;
sine[26571]=-65;
sine[26572]=-65;
sine[26573]=-65;
sine[26574]=-65;
sine[26575]=-65;
sine[26576]=-65;
sine[26577]=-65;
sine[26578]=-65;
sine[26579]=-65;
sine[26580]=-65;
sine[26581]=-65;
sine[26582]=-65;
sine[26583]=-66;
sine[26584]=-66;
sine[26585]=-66;
sine[26586]=-66;
sine[26587]=-66;
sine[26588]=-66;
sine[26589]=-66;
sine[26590]=-66;
sine[26591]=-66;
sine[26592]=-66;
sine[26593]=-66;
sine[26594]=-66;
sine[26595]=-66;
sine[26596]=-66;
sine[26597]=-66;
sine[26598]=-66;
sine[26599]=-66;
sine[26600]=-66;
sine[26601]=-66;
sine[26602]=-66;
sine[26603]=-66;
sine[26604]=-66;
sine[26605]=-66;
sine[26606]=-66;
sine[26607]=-66;
sine[26608]=-66;
sine[26609]=-66;
sine[26610]=-66;
sine[26611]=-66;
sine[26612]=-66;
sine[26613]=-66;
sine[26614]=-66;
sine[26615]=-66;
sine[26616]=-66;
sine[26617]=-66;
sine[26618]=-66;
sine[26619]=-66;
sine[26620]=-66;
sine[26621]=-67;
sine[26622]=-67;
sine[26623]=-67;
sine[26624]=-67;
sine[26625]=-67;
sine[26626]=-67;
sine[26627]=-67;
sine[26628]=-67;
sine[26629]=-67;
sine[26630]=-67;
sine[26631]=-67;
sine[26632]=-67;
sine[26633]=-67;
sine[26634]=-67;
sine[26635]=-67;
sine[26636]=-67;
sine[26637]=-67;
sine[26638]=-67;
sine[26639]=-67;
sine[26640]=-67;
sine[26641]=-67;
sine[26642]=-67;
sine[26643]=-67;
sine[26644]=-67;
sine[26645]=-67;
sine[26646]=-67;
sine[26647]=-67;
sine[26648]=-67;
sine[26649]=-67;
sine[26650]=-67;
sine[26651]=-67;
sine[26652]=-67;
sine[26653]=-67;
sine[26654]=-67;
sine[26655]=-67;
sine[26656]=-67;
sine[26657]=-67;
sine[26658]=-67;
sine[26659]=-67;
sine[26660]=-67;
sine[26661]=-68;
sine[26662]=-68;
sine[26663]=-68;
sine[26664]=-68;
sine[26665]=-68;
sine[26666]=-68;
sine[26667]=-68;
sine[26668]=-68;
sine[26669]=-68;
sine[26670]=-68;
sine[26671]=-68;
sine[26672]=-68;
sine[26673]=-68;
sine[26674]=-68;
sine[26675]=-68;
sine[26676]=-68;
sine[26677]=-68;
sine[26678]=-68;
sine[26679]=-68;
sine[26680]=-68;
sine[26681]=-68;
sine[26682]=-68;
sine[26683]=-68;
sine[26684]=-68;
sine[26685]=-68;
sine[26686]=-68;
sine[26687]=-68;
sine[26688]=-68;
sine[26689]=-68;
sine[26690]=-68;
sine[26691]=-68;
sine[26692]=-68;
sine[26693]=-68;
sine[26694]=-68;
sine[26695]=-68;
sine[26696]=-68;
sine[26697]=-68;
sine[26698]=-68;
sine[26699]=-68;
sine[26700]=-68;
sine[26701]=-68;
sine[26702]=-69;
sine[26703]=-69;
sine[26704]=-69;
sine[26705]=-69;
sine[26706]=-69;
sine[26707]=-69;
sine[26708]=-69;
sine[26709]=-69;
sine[26710]=-69;
sine[26711]=-69;
sine[26712]=-69;
sine[26713]=-69;
sine[26714]=-69;
sine[26715]=-69;
sine[26716]=-69;
sine[26717]=-69;
sine[26718]=-69;
sine[26719]=-69;
sine[26720]=-69;
sine[26721]=-69;
sine[26722]=-69;
sine[26723]=-69;
sine[26724]=-69;
sine[26725]=-69;
sine[26726]=-69;
sine[26727]=-69;
sine[26728]=-69;
sine[26729]=-69;
sine[26730]=-69;
sine[26731]=-69;
sine[26732]=-69;
sine[26733]=-69;
sine[26734]=-69;
sine[26735]=-69;
sine[26736]=-69;
sine[26737]=-69;
sine[26738]=-69;
sine[26739]=-69;
sine[26740]=-69;
sine[26741]=-69;
sine[26742]=-69;
sine[26743]=-69;
sine[26744]=-69;
sine[26745]=-69;
sine[26746]=-70;
sine[26747]=-70;
sine[26748]=-70;
sine[26749]=-70;
sine[26750]=-70;
sine[26751]=-70;
sine[26752]=-70;
sine[26753]=-70;
sine[26754]=-70;
sine[26755]=-70;
sine[26756]=-70;
sine[26757]=-70;
sine[26758]=-70;
sine[26759]=-70;
sine[26760]=-70;
sine[26761]=-70;
sine[26762]=-70;
sine[26763]=-70;
sine[26764]=-70;
sine[26765]=-70;
sine[26766]=-70;
sine[26767]=-70;
sine[26768]=-70;
sine[26769]=-70;
sine[26770]=-70;
sine[26771]=-70;
sine[26772]=-70;
sine[26773]=-70;
sine[26774]=-70;
sine[26775]=-70;
sine[26776]=-70;
sine[26777]=-70;
sine[26778]=-70;
sine[26779]=-70;
sine[26780]=-70;
sine[26781]=-70;
sine[26782]=-70;
sine[26783]=-70;
sine[26784]=-70;
sine[26785]=-70;
sine[26786]=-70;
sine[26787]=-70;
sine[26788]=-70;
sine[26789]=-70;
sine[26790]=-70;
sine[26791]=-71;
sine[26792]=-71;
sine[26793]=-71;
sine[26794]=-71;
sine[26795]=-71;
sine[26796]=-71;
sine[26797]=-71;
sine[26798]=-71;
sine[26799]=-71;
sine[26800]=-71;
sine[26801]=-71;
sine[26802]=-71;
sine[26803]=-71;
sine[26804]=-71;
sine[26805]=-71;
sine[26806]=-71;
sine[26807]=-71;
sine[26808]=-71;
sine[26809]=-71;
sine[26810]=-71;
sine[26811]=-71;
sine[26812]=-71;
sine[26813]=-71;
sine[26814]=-71;
sine[26815]=-71;
sine[26816]=-71;
sine[26817]=-71;
sine[26818]=-71;
sine[26819]=-71;
sine[26820]=-71;
sine[26821]=-71;
sine[26822]=-71;
sine[26823]=-71;
sine[26824]=-71;
sine[26825]=-71;
sine[26826]=-71;
sine[26827]=-71;
sine[26828]=-71;
sine[26829]=-71;
sine[26830]=-71;
sine[26831]=-71;
sine[26832]=-71;
sine[26833]=-71;
sine[26834]=-71;
sine[26835]=-71;
sine[26836]=-71;
sine[26837]=-71;
sine[26838]=-71;
sine[26839]=-71;
sine[26840]=-72;
sine[26841]=-72;
sine[26842]=-72;
sine[26843]=-72;
sine[26844]=-72;
sine[26845]=-72;
sine[26846]=-72;
sine[26847]=-72;
sine[26848]=-72;
sine[26849]=-72;
sine[26850]=-72;
sine[26851]=-72;
sine[26852]=-72;
sine[26853]=-72;
sine[26854]=-72;
sine[26855]=-72;
sine[26856]=-72;
sine[26857]=-72;
sine[26858]=-72;
sine[26859]=-72;
sine[26860]=-72;
sine[26861]=-72;
sine[26862]=-72;
sine[26863]=-72;
sine[26864]=-72;
sine[26865]=-72;
sine[26866]=-72;
sine[26867]=-72;
sine[26868]=-72;
sine[26869]=-72;
sine[26870]=-72;
sine[26871]=-72;
sine[26872]=-72;
sine[26873]=-72;
sine[26874]=-72;
sine[26875]=-72;
sine[26876]=-72;
sine[26877]=-72;
sine[26878]=-72;
sine[26879]=-72;
sine[26880]=-72;
sine[26881]=-72;
sine[26882]=-72;
sine[26883]=-72;
sine[26884]=-72;
sine[26885]=-72;
sine[26886]=-72;
sine[26887]=-72;
sine[26888]=-72;
sine[26889]=-72;
sine[26890]=-72;
sine[26891]=-72;
sine[26892]=-72;
sine[26893]=-73;
sine[26894]=-73;
sine[26895]=-73;
sine[26896]=-73;
sine[26897]=-73;
sine[26898]=-73;
sine[26899]=-73;
sine[26900]=-73;
sine[26901]=-73;
sine[26902]=-73;
sine[26903]=-73;
sine[26904]=-73;
sine[26905]=-73;
sine[26906]=-73;
sine[26907]=-73;
sine[26908]=-73;
sine[26909]=-73;
sine[26910]=-73;
sine[26911]=-73;
sine[26912]=-73;
sine[26913]=-73;
sine[26914]=-73;
sine[26915]=-73;
sine[26916]=-73;
sine[26917]=-73;
sine[26918]=-73;
sine[26919]=-73;
sine[26920]=-73;
sine[26921]=-73;
sine[26922]=-73;
sine[26923]=-73;
sine[26924]=-73;
sine[26925]=-73;
sine[26926]=-73;
sine[26927]=-73;
sine[26928]=-73;
sine[26929]=-73;
sine[26930]=-73;
sine[26931]=-73;
sine[26932]=-73;
sine[26933]=-73;
sine[26934]=-73;
sine[26935]=-73;
sine[26936]=-73;
sine[26937]=-73;
sine[26938]=-73;
sine[26939]=-73;
sine[26940]=-73;
sine[26941]=-73;
sine[26942]=-73;
sine[26943]=-73;
sine[26944]=-73;
sine[26945]=-73;
sine[26946]=-73;
sine[26947]=-73;
sine[26948]=-73;
sine[26949]=-73;
sine[26950]=-74;
sine[26951]=-74;
sine[26952]=-74;
sine[26953]=-74;
sine[26954]=-74;
sine[26955]=-74;
sine[26956]=-74;
sine[26957]=-74;
sine[26958]=-74;
sine[26959]=-74;
sine[26960]=-74;
sine[26961]=-74;
sine[26962]=-74;
sine[26963]=-74;
sine[26964]=-74;
sine[26965]=-74;
sine[26966]=-74;
sine[26967]=-74;
sine[26968]=-74;
sine[26969]=-74;
sine[26970]=-74;
sine[26971]=-74;
sine[26972]=-74;
sine[26973]=-74;
sine[26974]=-74;
sine[26975]=-74;
sine[26976]=-74;
sine[26977]=-74;
sine[26978]=-74;
sine[26979]=-74;
sine[26980]=-74;
sine[26981]=-74;
sine[26982]=-74;
sine[26983]=-74;
sine[26984]=-74;
sine[26985]=-74;
sine[26986]=-74;
sine[26987]=-74;
sine[26988]=-74;
sine[26989]=-74;
sine[26990]=-74;
sine[26991]=-74;
sine[26992]=-74;
sine[26993]=-74;
sine[26994]=-74;
sine[26995]=-74;
sine[26996]=-74;
sine[26997]=-74;
sine[26998]=-74;
sine[26999]=-74;
sine[27000]=-74;
sine[27001]=-74;
sine[27002]=-74;
sine[27003]=-74;
sine[27004]=-74;
sine[27005]=-74;
sine[27006]=-74;
sine[27007]=-74;
sine[27008]=-74;
sine[27009]=-74;
sine[27010]=-74;
sine[27011]=-74;
sine[27012]=-74;
sine[27013]=-74;
sine[27014]=-75;
sine[27015]=-75;
sine[27016]=-75;
sine[27017]=-75;
sine[27018]=-75;
sine[27019]=-75;
sine[27020]=-75;
sine[27021]=-75;
sine[27022]=-75;
sine[27023]=-75;
sine[27024]=-75;
sine[27025]=-75;
sine[27026]=-75;
sine[27027]=-75;
sine[27028]=-75;
sine[27029]=-75;
sine[27030]=-75;
sine[27031]=-75;
sine[27032]=-75;
sine[27033]=-75;
sine[27034]=-75;
sine[27035]=-75;
sine[27036]=-75;
sine[27037]=-75;
sine[27038]=-75;
sine[27039]=-75;
sine[27040]=-75;
sine[27041]=-75;
sine[27042]=-75;
sine[27043]=-75;
sine[27044]=-75;
sine[27045]=-75;
sine[27046]=-75;
sine[27047]=-75;
sine[27048]=-75;
sine[27049]=-75;
sine[27050]=-75;
sine[27051]=-75;
sine[27052]=-75;
sine[27053]=-75;
sine[27054]=-75;
sine[27055]=-75;
sine[27056]=-75;
sine[27057]=-75;
sine[27058]=-75;
sine[27059]=-75;
sine[27060]=-75;
sine[27061]=-75;
sine[27062]=-75;
sine[27063]=-75;
sine[27064]=-75;
sine[27065]=-75;
sine[27066]=-75;
sine[27067]=-75;
sine[27068]=-75;
sine[27069]=-75;
sine[27070]=-75;
sine[27071]=-75;
sine[27072]=-75;
sine[27073]=-75;
sine[27074]=-75;
sine[27075]=-75;
sine[27076]=-75;
sine[27077]=-75;
sine[27078]=-75;
sine[27079]=-75;
sine[27080]=-75;
sine[27081]=-75;
sine[27082]=-75;
sine[27083]=-75;
sine[27084]=-75;
sine[27085]=-75;
sine[27086]=-75;
sine[27087]=-76;
sine[27088]=-76;
sine[27089]=-76;
sine[27090]=-76;
sine[27091]=-76;
sine[27092]=-76;
sine[27093]=-76;
sine[27094]=-76;
sine[27095]=-76;
sine[27096]=-76;
sine[27097]=-76;
sine[27098]=-76;
sine[27099]=-76;
sine[27100]=-76;
sine[27101]=-76;
sine[27102]=-76;
sine[27103]=-76;
sine[27104]=-76;
sine[27105]=-76;
sine[27106]=-76;
sine[27107]=-76;
sine[27108]=-76;
sine[27109]=-76;
sine[27110]=-76;
sine[27111]=-76;
sine[27112]=-76;
sine[27113]=-76;
sine[27114]=-76;
sine[27115]=-76;
sine[27116]=-76;
sine[27117]=-76;
sine[27118]=-76;
sine[27119]=-76;
sine[27120]=-76;
sine[27121]=-76;
sine[27122]=-76;
sine[27123]=-76;
sine[27124]=-76;
sine[27125]=-76;
sine[27126]=-76;
sine[27127]=-76;
sine[27128]=-76;
sine[27129]=-76;
sine[27130]=-76;
sine[27131]=-76;
sine[27132]=-76;
sine[27133]=-76;
sine[27134]=-76;
sine[27135]=-76;
sine[27136]=-76;
sine[27137]=-76;
sine[27138]=-76;
sine[27139]=-76;
sine[27140]=-76;
sine[27141]=-76;
sine[27142]=-76;
sine[27143]=-76;
sine[27144]=-76;
sine[27145]=-76;
sine[27146]=-76;
sine[27147]=-76;
sine[27148]=-76;
sine[27149]=-76;
sine[27150]=-76;
sine[27151]=-76;
sine[27152]=-76;
sine[27153]=-76;
sine[27154]=-76;
sine[27155]=-76;
sine[27156]=-76;
sine[27157]=-76;
sine[27158]=-76;
sine[27159]=-76;
sine[27160]=-76;
sine[27161]=-76;
sine[27162]=-76;
sine[27163]=-76;
sine[27164]=-76;
sine[27165]=-76;
sine[27166]=-76;
sine[27167]=-76;
sine[27168]=-76;
sine[27169]=-76;
sine[27170]=-76;
sine[27171]=-76;
sine[27172]=-76;
sine[27173]=-76;
sine[27174]=-76;
sine[27175]=-77;
sine[27176]=-77;
sine[27177]=-77;
sine[27178]=-77;
sine[27179]=-77;
sine[27180]=-77;
sine[27181]=-77;
sine[27182]=-77;
sine[27183]=-77;
sine[27184]=-77;
sine[27185]=-77;
sine[27186]=-77;
sine[27187]=-77;
sine[27188]=-77;
sine[27189]=-77;
sine[27190]=-77;
sine[27191]=-77;
sine[27192]=-77;
sine[27193]=-77;
sine[27194]=-77;
sine[27195]=-77;
sine[27196]=-77;
sine[27197]=-77;
sine[27198]=-77;
sine[27199]=-77;
sine[27200]=-77;
sine[27201]=-77;
sine[27202]=-77;
sine[27203]=-77;
sine[27204]=-77;
sine[27205]=-77;
sine[27206]=-77;
sine[27207]=-77;
sine[27208]=-77;
sine[27209]=-77;
sine[27210]=-77;
sine[27211]=-77;
sine[27212]=-77;
sine[27213]=-77;
sine[27214]=-77;
sine[27215]=-77;
sine[27216]=-77;
sine[27217]=-77;
sine[27218]=-77;
sine[27219]=-77;
sine[27220]=-77;
sine[27221]=-77;
sine[27222]=-77;
sine[27223]=-77;
sine[27224]=-77;
sine[27225]=-77;
sine[27226]=-77;
sine[27227]=-77;
sine[27228]=-77;
sine[27229]=-77;
sine[27230]=-77;
sine[27231]=-77;
sine[27232]=-77;
sine[27233]=-77;
sine[27234]=-77;
sine[27235]=-77;
sine[27236]=-77;
sine[27237]=-77;
sine[27238]=-77;
sine[27239]=-77;
sine[27240]=-77;
sine[27241]=-77;
sine[27242]=-77;
sine[27243]=-77;
sine[27244]=-77;
sine[27245]=-77;
sine[27246]=-77;
sine[27247]=-77;
sine[27248]=-77;
sine[27249]=-77;
sine[27250]=-77;
sine[27251]=-77;
sine[27252]=-77;
sine[27253]=-77;
sine[27254]=-77;
sine[27255]=-77;
sine[27256]=-77;
sine[27257]=-77;
sine[27258]=-77;
sine[27259]=-77;
sine[27260]=-77;
sine[27261]=-77;
sine[27262]=-77;
sine[27263]=-77;
sine[27264]=-77;
sine[27265]=-77;
sine[27266]=-77;
sine[27267]=-77;
sine[27268]=-77;
sine[27269]=-77;
sine[27270]=-77;
sine[27271]=-77;
sine[27272]=-77;
sine[27273]=-77;
sine[27274]=-77;
sine[27275]=-77;
sine[27276]=-77;
sine[27277]=-77;
sine[27278]=-77;
sine[27279]=-77;
sine[27280]=-77;
sine[27281]=-77;
sine[27282]=-77;
sine[27283]=-77;
sine[27284]=-77;
sine[27285]=-77;
sine[27286]=-77;
sine[27287]=-77;
sine[27288]=-77;
sine[27289]=-77;
sine[27290]=-77;
sine[27291]=-77;
sine[27292]=-77;
sine[27293]=-77;
sine[27294]=-77;
sine[27295]=-77;
sine[27296]=-77;
sine[27297]=-77;
sine[27298]=-77;
sine[27299]=-78;
sine[27300]=-78;
sine[27301]=-78;
sine[27302]=-78;
sine[27303]=-78;
sine[27304]=-78;
sine[27305]=-78;
sine[27306]=-78;
sine[27307]=-78;
sine[27308]=-78;
sine[27309]=-78;
sine[27310]=-78;
sine[27311]=-78;
sine[27312]=-78;
sine[27313]=-78;
sine[27314]=-78;
sine[27315]=-78;
sine[27316]=-78;
sine[27317]=-78;
sine[27318]=-78;
sine[27319]=-78;
sine[27320]=-78;
sine[27321]=-78;
sine[27322]=-78;
sine[27323]=-78;
sine[27324]=-78;
sine[27325]=-78;
sine[27326]=-78;
sine[27327]=-78;
sine[27328]=-78;
sine[27329]=-78;
sine[27330]=-78;
sine[27331]=-78;
sine[27332]=-78;
sine[27333]=-78;
sine[27334]=-78;
sine[27335]=-78;
sine[27336]=-78;
sine[27337]=-78;
sine[27338]=-78;
sine[27339]=-78;
sine[27340]=-78;
sine[27341]=-78;
sine[27342]=-78;
sine[27343]=-78;
sine[27344]=-78;
sine[27345]=-78;
sine[27346]=-78;
sine[27347]=-78;
sine[27348]=-78;
sine[27349]=-78;
sine[27350]=-78;
sine[27351]=-78;
sine[27352]=-78;
sine[27353]=-78;
sine[27354]=-78;
sine[27355]=-78;
sine[27356]=-78;
sine[27357]=-78;
sine[27358]=-78;
sine[27359]=-78;
sine[27360]=-78;
sine[27361]=-78;
sine[27362]=-78;
sine[27363]=-78;
sine[27364]=-78;
sine[27365]=-78;
sine[27366]=-78;
sine[27367]=-78;
sine[27368]=-78;
sine[27369]=-78;
sine[27370]=-78;
sine[27371]=-78;
sine[27372]=-78;
sine[27373]=-78;
sine[27374]=-78;
sine[27375]=-78;
sine[27376]=-78;
sine[27377]=-78;
sine[27378]=-78;
sine[27379]=-78;
sine[27380]=-78;
sine[27381]=-78;
sine[27382]=-78;
sine[27383]=-78;
sine[27384]=-78;
sine[27385]=-78;
sine[27386]=-78;
sine[27387]=-78;
sine[27388]=-78;
sine[27389]=-78;
sine[27390]=-78;
sine[27391]=-78;
sine[27392]=-78;
sine[27393]=-78;
sine[27394]=-78;
sine[27395]=-78;
sine[27396]=-78;
sine[27397]=-78;
sine[27398]=-78;
sine[27399]=-78;
sine[27400]=-78;
sine[27401]=-78;
sine[27402]=-78;
sine[27403]=-78;
sine[27404]=-78;
sine[27405]=-78;
sine[27406]=-78;
sine[27407]=-78;
sine[27408]=-78;
sine[27409]=-78;
sine[27410]=-78;
sine[27411]=-78;
sine[27412]=-78;
sine[27413]=-78;
sine[27414]=-78;
sine[27415]=-78;
sine[27416]=-78;
sine[27417]=-78;
sine[27418]=-78;
sine[27419]=-78;
sine[27420]=-78;
sine[27421]=-78;
sine[27422]=-78;
sine[27423]=-78;
sine[27424]=-78;
sine[27425]=-78;
sine[27426]=-78;
sine[27427]=-78;
sine[27428]=-78;
sine[27429]=-78;
sine[27430]=-78;
sine[27431]=-78;
sine[27432]=-78;
sine[27433]=-78;
sine[27434]=-78;
sine[27435]=-78;
sine[27436]=-78;
sine[27437]=-78;
sine[27438]=-78;
sine[27439]=-78;
sine[27440]=-78;
sine[27441]=-78;
sine[27442]=-78;
sine[27443]=-78;
sine[27444]=-78;
sine[27445]=-78;
sine[27446]=-78;
sine[27447]=-78;
sine[27448]=-78;
sine[27449]=-78;
sine[27450]=-78;
sine[27451]=-78;
sine[27452]=-78;
sine[27453]=-78;
sine[27454]=-78;
sine[27455]=-78;
sine[27456]=-78;
sine[27457]=-78;
sine[27458]=-78;
sine[27459]=-78;
sine[27460]=-78;
sine[27461]=-78;
sine[27462]=-78;
sine[27463]=-78;
sine[27464]=-78;
sine[27465]=-78;
sine[27466]=-78;
sine[27467]=-78;
sine[27468]=-78;
sine[27469]=-78;
sine[27470]=-78;
sine[27471]=-78;
sine[27472]=-78;
sine[27473]=-78;
sine[27474]=-78;
sine[27475]=-78;
sine[27476]=-78;
sine[27477]=-78;
sine[27478]=-78;
sine[27479]=-78;
sine[27480]=-78;
sine[27481]=-78;
sine[27482]=-78;
sine[27483]=-78;
sine[27484]=-78;
sine[27485]=-78;
sine[27486]=-78;
sine[27487]=-78;
sine[27488]=-78;
sine[27489]=-78;
sine[27490]=-78;
sine[27491]=-78;
sine[27492]=-78;
sine[27493]=-78;
sine[27494]=-78;
sine[27495]=-78;
sine[27496]=-78;
sine[27497]=-78;
sine[27498]=-78;
sine[27499]=-78;
sine[27500]=-78;
sine[27501]=-78;
sine[27502]=-78;
sine[27503]=-78;
sine[27504]=-78;
sine[27505]=-78;
sine[27506]=-78;
sine[27507]=-78;
sine[27508]=-78;
sine[27509]=-78;
sine[27510]=-78;
sine[27511]=-78;
sine[27512]=-78;
sine[27513]=-78;
sine[27514]=-78;
sine[27515]=-78;
sine[27516]=-78;
sine[27517]=-78;
sine[27518]=-78;
sine[27519]=-78;
sine[27520]=-78;
sine[27521]=-78;
sine[27522]=-78;
sine[27523]=-78;
sine[27524]=-78;
sine[27525]=-78;
sine[27526]=-78;
sine[27527]=-78;
sine[27528]=-78;
sine[27529]=-78;
sine[27530]=-78;
sine[27531]=-78;
sine[27532]=-78;
sine[27533]=-78;
sine[27534]=-78;
sine[27535]=-78;
sine[27536]=-78;
sine[27537]=-78;
sine[27538]=-78;
sine[27539]=-78;
sine[27540]=-78;
sine[27541]=-78;
sine[27542]=-78;
sine[27543]=-78;
sine[27544]=-78;
sine[27545]=-78;
sine[27546]=-78;
sine[27547]=-78;
sine[27548]=-78;
sine[27549]=-78;
sine[27550]=-78;
sine[27551]=-78;
sine[27552]=-78;
sine[27553]=-78;
sine[27554]=-78;
sine[27555]=-78;
sine[27556]=-78;
sine[27557]=-78;
sine[27558]=-78;
sine[27559]=-78;
sine[27560]=-78;
sine[27561]=-78;
sine[27562]=-78;
sine[27563]=-78;
sine[27564]=-78;
sine[27565]=-78;
sine[27566]=-78;
sine[27567]=-78;
sine[27568]=-78;
sine[27569]=-78;
sine[27570]=-78;
sine[27571]=-78;
sine[27572]=-78;
sine[27573]=-78;
sine[27574]=-78;
sine[27575]=-78;
sine[27576]=-78;
sine[27577]=-78;
sine[27578]=-78;
sine[27579]=-78;
sine[27580]=-78;
sine[27581]=-78;
sine[27582]=-78;
sine[27583]=-78;
sine[27584]=-78;
sine[27585]=-78;
sine[27586]=-78;
sine[27587]=-78;
sine[27588]=-78;
sine[27589]=-78;
sine[27590]=-78;
sine[27591]=-78;
sine[27592]=-78;
sine[27593]=-78;
sine[27594]=-78;
sine[27595]=-78;
sine[27596]=-78;
sine[27597]=-78;
sine[27598]=-78;
sine[27599]=-78;
sine[27600]=-78;
sine[27601]=-78;
sine[27602]=-78;
sine[27603]=-78;
sine[27604]=-78;
sine[27605]=-78;
sine[27606]=-78;
sine[27607]=-78;
sine[27608]=-78;
sine[27609]=-78;
sine[27610]=-78;
sine[27611]=-78;
sine[27612]=-78;
sine[27613]=-78;
sine[27614]=-78;
sine[27615]=-78;
sine[27616]=-78;
sine[27617]=-78;
sine[27618]=-78;
sine[27619]=-78;
sine[27620]=-78;
sine[27621]=-78;
sine[27622]=-78;
sine[27623]=-78;
sine[27624]=-78;
sine[27625]=-78;
sine[27626]=-78;
sine[27627]=-78;
sine[27628]=-78;
sine[27629]=-78;
sine[27630]=-78;
sine[27631]=-78;
sine[27632]=-78;
sine[27633]=-78;
sine[27634]=-78;
sine[27635]=-78;
sine[27636]=-78;
sine[27637]=-78;
sine[27638]=-78;
sine[27639]=-78;
sine[27640]=-78;
sine[27641]=-78;
sine[27642]=-78;
sine[27643]=-78;
sine[27644]=-78;
sine[27645]=-78;
sine[27646]=-78;
sine[27647]=-78;
sine[27648]=-78;
sine[27649]=-78;
sine[27650]=-78;
sine[27651]=-78;
sine[27652]=-78;
sine[27653]=-78;
sine[27654]=-78;
sine[27655]=-78;
sine[27656]=-78;
sine[27657]=-78;
sine[27658]=-78;
sine[27659]=-78;
sine[27660]=-78;
sine[27661]=-78;
sine[27662]=-78;
sine[27663]=-78;
sine[27664]=-78;
sine[27665]=-78;
sine[27666]=-78;
sine[27667]=-78;
sine[27668]=-78;
sine[27669]=-78;
sine[27670]=-78;
sine[27671]=-78;
sine[27672]=-78;
sine[27673]=-78;
sine[27674]=-78;
sine[27675]=-78;
sine[27676]=-78;
sine[27677]=-78;
sine[27678]=-78;
sine[27679]=-78;
sine[27680]=-78;
sine[27681]=-78;
sine[27682]=-78;
sine[27683]=-78;
sine[27684]=-78;
sine[27685]=-78;
sine[27686]=-78;
sine[27687]=-78;
sine[27688]=-78;
sine[27689]=-78;
sine[27690]=-78;
sine[27691]=-78;
sine[27692]=-78;
sine[27693]=-78;
sine[27694]=-78;
sine[27695]=-78;
sine[27696]=-78;
sine[27697]=-78;
sine[27698]=-78;
sine[27699]=-78;
sine[27700]=-78;
sine[27701]=-78;
sine[27702]=-77;
sine[27703]=-77;
sine[27704]=-77;
sine[27705]=-77;
sine[27706]=-77;
sine[27707]=-77;
sine[27708]=-77;
sine[27709]=-77;
sine[27710]=-77;
sine[27711]=-77;
sine[27712]=-77;
sine[27713]=-77;
sine[27714]=-77;
sine[27715]=-77;
sine[27716]=-77;
sine[27717]=-77;
sine[27718]=-77;
sine[27719]=-77;
sine[27720]=-77;
sine[27721]=-77;
sine[27722]=-77;
sine[27723]=-77;
sine[27724]=-77;
sine[27725]=-77;
sine[27726]=-77;
sine[27727]=-77;
sine[27728]=-77;
sine[27729]=-77;
sine[27730]=-77;
sine[27731]=-77;
sine[27732]=-77;
sine[27733]=-77;
sine[27734]=-77;
sine[27735]=-77;
sine[27736]=-77;
sine[27737]=-77;
sine[27738]=-77;
sine[27739]=-77;
sine[27740]=-77;
sine[27741]=-77;
sine[27742]=-77;
sine[27743]=-77;
sine[27744]=-77;
sine[27745]=-77;
sine[27746]=-77;
sine[27747]=-77;
sine[27748]=-77;
sine[27749]=-77;
sine[27750]=-77;
sine[27751]=-77;
sine[27752]=-77;
sine[27753]=-77;
sine[27754]=-77;
sine[27755]=-77;
sine[27756]=-77;
sine[27757]=-77;
sine[27758]=-77;
sine[27759]=-77;
sine[27760]=-77;
sine[27761]=-77;
sine[27762]=-77;
sine[27763]=-77;
sine[27764]=-77;
sine[27765]=-77;
sine[27766]=-77;
sine[27767]=-77;
sine[27768]=-77;
sine[27769]=-77;
sine[27770]=-77;
sine[27771]=-77;
sine[27772]=-77;
sine[27773]=-77;
sine[27774]=-77;
sine[27775]=-77;
sine[27776]=-77;
sine[27777]=-77;
sine[27778]=-77;
sine[27779]=-77;
sine[27780]=-77;
sine[27781]=-77;
sine[27782]=-77;
sine[27783]=-77;
sine[27784]=-77;
sine[27785]=-77;
sine[27786]=-77;
sine[27787]=-77;
sine[27788]=-77;
sine[27789]=-77;
sine[27790]=-77;
sine[27791]=-77;
sine[27792]=-77;
sine[27793]=-77;
sine[27794]=-77;
sine[27795]=-77;
sine[27796]=-77;
sine[27797]=-77;
sine[27798]=-77;
sine[27799]=-77;
sine[27800]=-77;
sine[27801]=-77;
sine[27802]=-77;
sine[27803]=-77;
sine[27804]=-77;
sine[27805]=-77;
sine[27806]=-77;
sine[27807]=-77;
sine[27808]=-77;
sine[27809]=-77;
sine[27810]=-77;
sine[27811]=-77;
sine[27812]=-77;
sine[27813]=-77;
sine[27814]=-77;
sine[27815]=-77;
sine[27816]=-77;
sine[27817]=-77;
sine[27818]=-77;
sine[27819]=-77;
sine[27820]=-77;
sine[27821]=-77;
sine[27822]=-77;
sine[27823]=-77;
sine[27824]=-77;
sine[27825]=-77;
sine[27826]=-76;
sine[27827]=-76;
sine[27828]=-76;
sine[27829]=-76;
sine[27830]=-76;
sine[27831]=-76;
sine[27832]=-76;
sine[27833]=-76;
sine[27834]=-76;
sine[27835]=-76;
sine[27836]=-76;
sine[27837]=-76;
sine[27838]=-76;
sine[27839]=-76;
sine[27840]=-76;
sine[27841]=-76;
sine[27842]=-76;
sine[27843]=-76;
sine[27844]=-76;
sine[27845]=-76;
sine[27846]=-76;
sine[27847]=-76;
sine[27848]=-76;
sine[27849]=-76;
sine[27850]=-76;
sine[27851]=-76;
sine[27852]=-76;
sine[27853]=-76;
sine[27854]=-76;
sine[27855]=-76;
sine[27856]=-76;
sine[27857]=-76;
sine[27858]=-76;
sine[27859]=-76;
sine[27860]=-76;
sine[27861]=-76;
sine[27862]=-76;
sine[27863]=-76;
sine[27864]=-76;
sine[27865]=-76;
sine[27866]=-76;
sine[27867]=-76;
sine[27868]=-76;
sine[27869]=-76;
sine[27870]=-76;
sine[27871]=-76;
sine[27872]=-76;
sine[27873]=-76;
sine[27874]=-76;
sine[27875]=-76;
sine[27876]=-76;
sine[27877]=-76;
sine[27878]=-76;
sine[27879]=-76;
sine[27880]=-76;
sine[27881]=-76;
sine[27882]=-76;
sine[27883]=-76;
sine[27884]=-76;
sine[27885]=-76;
sine[27886]=-76;
sine[27887]=-76;
sine[27888]=-76;
sine[27889]=-76;
sine[27890]=-76;
sine[27891]=-76;
sine[27892]=-76;
sine[27893]=-76;
sine[27894]=-76;
sine[27895]=-76;
sine[27896]=-76;
sine[27897]=-76;
sine[27898]=-76;
sine[27899]=-76;
sine[27900]=-76;
sine[27901]=-76;
sine[27902]=-76;
sine[27903]=-76;
sine[27904]=-76;
sine[27905]=-76;
sine[27906]=-76;
sine[27907]=-76;
sine[27908]=-76;
sine[27909]=-76;
sine[27910]=-76;
sine[27911]=-76;
sine[27912]=-76;
sine[27913]=-76;
sine[27914]=-75;
sine[27915]=-75;
sine[27916]=-75;
sine[27917]=-75;
sine[27918]=-75;
sine[27919]=-75;
sine[27920]=-75;
sine[27921]=-75;
sine[27922]=-75;
sine[27923]=-75;
sine[27924]=-75;
sine[27925]=-75;
sine[27926]=-75;
sine[27927]=-75;
sine[27928]=-75;
sine[27929]=-75;
sine[27930]=-75;
sine[27931]=-75;
sine[27932]=-75;
sine[27933]=-75;
sine[27934]=-75;
sine[27935]=-75;
sine[27936]=-75;
sine[27937]=-75;
sine[27938]=-75;
sine[27939]=-75;
sine[27940]=-75;
sine[27941]=-75;
sine[27942]=-75;
sine[27943]=-75;
sine[27944]=-75;
sine[27945]=-75;
sine[27946]=-75;
sine[27947]=-75;
sine[27948]=-75;
sine[27949]=-75;
sine[27950]=-75;
sine[27951]=-75;
sine[27952]=-75;
sine[27953]=-75;
sine[27954]=-75;
sine[27955]=-75;
sine[27956]=-75;
sine[27957]=-75;
sine[27958]=-75;
sine[27959]=-75;
sine[27960]=-75;
sine[27961]=-75;
sine[27962]=-75;
sine[27963]=-75;
sine[27964]=-75;
sine[27965]=-75;
sine[27966]=-75;
sine[27967]=-75;
sine[27968]=-75;
sine[27969]=-75;
sine[27970]=-75;
sine[27971]=-75;
sine[27972]=-75;
sine[27973]=-75;
sine[27974]=-75;
sine[27975]=-75;
sine[27976]=-75;
sine[27977]=-75;
sine[27978]=-75;
sine[27979]=-75;
sine[27980]=-75;
sine[27981]=-75;
sine[27982]=-75;
sine[27983]=-75;
sine[27984]=-75;
sine[27985]=-75;
sine[27986]=-75;
sine[27987]=-74;
sine[27988]=-74;
sine[27989]=-74;
sine[27990]=-74;
sine[27991]=-74;
sine[27992]=-74;
sine[27993]=-74;
sine[27994]=-74;
sine[27995]=-74;
sine[27996]=-74;
sine[27997]=-74;
sine[27998]=-74;
sine[27999]=-74;
sine[28000]=-74;
sine[28001]=-74;
sine[28002]=-74;
sine[28003]=-74;
sine[28004]=-74;
sine[28005]=-74;
sine[28006]=-74;
sine[28007]=-74;
sine[28008]=-74;
sine[28009]=-74;
sine[28010]=-74;
sine[28011]=-74;
sine[28012]=-74;
sine[28013]=-74;
sine[28014]=-74;
sine[28015]=-74;
sine[28016]=-74;
sine[28017]=-74;
sine[28018]=-74;
sine[28019]=-74;
sine[28020]=-74;
sine[28021]=-74;
sine[28022]=-74;
sine[28023]=-74;
sine[28024]=-74;
sine[28025]=-74;
sine[28026]=-74;
sine[28027]=-74;
sine[28028]=-74;
sine[28029]=-74;
sine[28030]=-74;
sine[28031]=-74;
sine[28032]=-74;
sine[28033]=-74;
sine[28034]=-74;
sine[28035]=-74;
sine[28036]=-74;
sine[28037]=-74;
sine[28038]=-74;
sine[28039]=-74;
sine[28040]=-74;
sine[28041]=-74;
sine[28042]=-74;
sine[28043]=-74;
sine[28044]=-74;
sine[28045]=-74;
sine[28046]=-74;
sine[28047]=-74;
sine[28048]=-74;
sine[28049]=-74;
sine[28050]=-74;
sine[28051]=-73;
sine[28052]=-73;
sine[28053]=-73;
sine[28054]=-73;
sine[28055]=-73;
sine[28056]=-73;
sine[28057]=-73;
sine[28058]=-73;
sine[28059]=-73;
sine[28060]=-73;
sine[28061]=-73;
sine[28062]=-73;
sine[28063]=-73;
sine[28064]=-73;
sine[28065]=-73;
sine[28066]=-73;
sine[28067]=-73;
sine[28068]=-73;
sine[28069]=-73;
sine[28070]=-73;
sine[28071]=-73;
sine[28072]=-73;
sine[28073]=-73;
sine[28074]=-73;
sine[28075]=-73;
sine[28076]=-73;
sine[28077]=-73;
sine[28078]=-73;
sine[28079]=-73;
sine[28080]=-73;
sine[28081]=-73;
sine[28082]=-73;
sine[28083]=-73;
sine[28084]=-73;
sine[28085]=-73;
sine[28086]=-73;
sine[28087]=-73;
sine[28088]=-73;
sine[28089]=-73;
sine[28090]=-73;
sine[28091]=-73;
sine[28092]=-73;
sine[28093]=-73;
sine[28094]=-73;
sine[28095]=-73;
sine[28096]=-73;
sine[28097]=-73;
sine[28098]=-73;
sine[28099]=-73;
sine[28100]=-73;
sine[28101]=-73;
sine[28102]=-73;
sine[28103]=-73;
sine[28104]=-73;
sine[28105]=-73;
sine[28106]=-73;
sine[28107]=-73;
sine[28108]=-72;
sine[28109]=-72;
sine[28110]=-72;
sine[28111]=-72;
sine[28112]=-72;
sine[28113]=-72;
sine[28114]=-72;
sine[28115]=-72;
sine[28116]=-72;
sine[28117]=-72;
sine[28118]=-72;
sine[28119]=-72;
sine[28120]=-72;
sine[28121]=-72;
sine[28122]=-72;
sine[28123]=-72;
sine[28124]=-72;
sine[28125]=-72;
sine[28126]=-72;
sine[28127]=-72;
sine[28128]=-72;
sine[28129]=-72;
sine[28130]=-72;
sine[28131]=-72;
sine[28132]=-72;
sine[28133]=-72;
sine[28134]=-72;
sine[28135]=-72;
sine[28136]=-72;
sine[28137]=-72;
sine[28138]=-72;
sine[28139]=-72;
sine[28140]=-72;
sine[28141]=-72;
sine[28142]=-72;
sine[28143]=-72;
sine[28144]=-72;
sine[28145]=-72;
sine[28146]=-72;
sine[28147]=-72;
sine[28148]=-72;
sine[28149]=-72;
sine[28150]=-72;
sine[28151]=-72;
sine[28152]=-72;
sine[28153]=-72;
sine[28154]=-72;
sine[28155]=-72;
sine[28156]=-72;
sine[28157]=-72;
sine[28158]=-72;
sine[28159]=-72;
sine[28160]=-72;
sine[28161]=-71;
sine[28162]=-71;
sine[28163]=-71;
sine[28164]=-71;
sine[28165]=-71;
sine[28166]=-71;
sine[28167]=-71;
sine[28168]=-71;
sine[28169]=-71;
sine[28170]=-71;
sine[28171]=-71;
sine[28172]=-71;
sine[28173]=-71;
sine[28174]=-71;
sine[28175]=-71;
sine[28176]=-71;
sine[28177]=-71;
sine[28178]=-71;
sine[28179]=-71;
sine[28180]=-71;
sine[28181]=-71;
sine[28182]=-71;
sine[28183]=-71;
sine[28184]=-71;
sine[28185]=-71;
sine[28186]=-71;
sine[28187]=-71;
sine[28188]=-71;
sine[28189]=-71;
sine[28190]=-71;
sine[28191]=-71;
sine[28192]=-71;
sine[28193]=-71;
sine[28194]=-71;
sine[28195]=-71;
sine[28196]=-71;
sine[28197]=-71;
sine[28198]=-71;
sine[28199]=-71;
sine[28200]=-71;
sine[28201]=-71;
sine[28202]=-71;
sine[28203]=-71;
sine[28204]=-71;
sine[28205]=-71;
sine[28206]=-71;
sine[28207]=-71;
sine[28208]=-71;
sine[28209]=-71;
sine[28210]=-70;
sine[28211]=-70;
sine[28212]=-70;
sine[28213]=-70;
sine[28214]=-70;
sine[28215]=-70;
sine[28216]=-70;
sine[28217]=-70;
sine[28218]=-70;
sine[28219]=-70;
sine[28220]=-70;
sine[28221]=-70;
sine[28222]=-70;
sine[28223]=-70;
sine[28224]=-70;
sine[28225]=-70;
sine[28226]=-70;
sine[28227]=-70;
sine[28228]=-70;
sine[28229]=-70;
sine[28230]=-70;
sine[28231]=-70;
sine[28232]=-70;
sine[28233]=-70;
sine[28234]=-70;
sine[28235]=-70;
sine[28236]=-70;
sine[28237]=-70;
sine[28238]=-70;
sine[28239]=-70;
sine[28240]=-70;
sine[28241]=-70;
sine[28242]=-70;
sine[28243]=-70;
sine[28244]=-70;
sine[28245]=-70;
sine[28246]=-70;
sine[28247]=-70;
sine[28248]=-70;
sine[28249]=-70;
sine[28250]=-70;
sine[28251]=-70;
sine[28252]=-70;
sine[28253]=-70;
sine[28254]=-70;
sine[28255]=-69;
sine[28256]=-69;
sine[28257]=-69;
sine[28258]=-69;
sine[28259]=-69;
sine[28260]=-69;
sine[28261]=-69;
sine[28262]=-69;
sine[28263]=-69;
sine[28264]=-69;
sine[28265]=-69;
sine[28266]=-69;
sine[28267]=-69;
sine[28268]=-69;
sine[28269]=-69;
sine[28270]=-69;
sine[28271]=-69;
sine[28272]=-69;
sine[28273]=-69;
sine[28274]=-69;
sine[28275]=-69;
sine[28276]=-69;
sine[28277]=-69;
sine[28278]=-69;
sine[28279]=-69;
sine[28280]=-69;
sine[28281]=-69;
sine[28282]=-69;
sine[28283]=-69;
sine[28284]=-69;
sine[28285]=-69;
sine[28286]=-69;
sine[28287]=-69;
sine[28288]=-69;
sine[28289]=-69;
sine[28290]=-69;
sine[28291]=-69;
sine[28292]=-69;
sine[28293]=-69;
sine[28294]=-69;
sine[28295]=-69;
sine[28296]=-69;
sine[28297]=-69;
sine[28298]=-69;
sine[28299]=-68;
sine[28300]=-68;
sine[28301]=-68;
sine[28302]=-68;
sine[28303]=-68;
sine[28304]=-68;
sine[28305]=-68;
sine[28306]=-68;
sine[28307]=-68;
sine[28308]=-68;
sine[28309]=-68;
sine[28310]=-68;
sine[28311]=-68;
sine[28312]=-68;
sine[28313]=-68;
sine[28314]=-68;
sine[28315]=-68;
sine[28316]=-68;
sine[28317]=-68;
sine[28318]=-68;
sine[28319]=-68;
sine[28320]=-68;
sine[28321]=-68;
sine[28322]=-68;
sine[28323]=-68;
sine[28324]=-68;
sine[28325]=-68;
sine[28326]=-68;
sine[28327]=-68;
sine[28328]=-68;
sine[28329]=-68;
sine[28330]=-68;
sine[28331]=-68;
sine[28332]=-68;
sine[28333]=-68;
sine[28334]=-68;
sine[28335]=-68;
sine[28336]=-68;
sine[28337]=-68;
sine[28338]=-68;
sine[28339]=-68;
sine[28340]=-67;
sine[28341]=-67;
sine[28342]=-67;
sine[28343]=-67;
sine[28344]=-67;
sine[28345]=-67;
sine[28346]=-67;
sine[28347]=-67;
sine[28348]=-67;
sine[28349]=-67;
sine[28350]=-67;
sine[28351]=-67;
sine[28352]=-67;
sine[28353]=-67;
sine[28354]=-67;
sine[28355]=-67;
sine[28356]=-67;
sine[28357]=-67;
sine[28358]=-67;
sine[28359]=-67;
sine[28360]=-67;
sine[28361]=-67;
sine[28362]=-67;
sine[28363]=-67;
sine[28364]=-67;
sine[28365]=-67;
sine[28366]=-67;
sine[28367]=-67;
sine[28368]=-67;
sine[28369]=-67;
sine[28370]=-67;
sine[28371]=-67;
sine[28372]=-67;
sine[28373]=-67;
sine[28374]=-67;
sine[28375]=-67;
sine[28376]=-67;
sine[28377]=-67;
sine[28378]=-67;
sine[28379]=-67;
sine[28380]=-66;
sine[28381]=-66;
sine[28382]=-66;
sine[28383]=-66;
sine[28384]=-66;
sine[28385]=-66;
sine[28386]=-66;
sine[28387]=-66;
sine[28388]=-66;
sine[28389]=-66;
sine[28390]=-66;
sine[28391]=-66;
sine[28392]=-66;
sine[28393]=-66;
sine[28394]=-66;
sine[28395]=-66;
sine[28396]=-66;
sine[28397]=-66;
sine[28398]=-66;
sine[28399]=-66;
sine[28400]=-66;
sine[28401]=-66;
sine[28402]=-66;
sine[28403]=-66;
sine[28404]=-66;
sine[28405]=-66;
sine[28406]=-66;
sine[28407]=-66;
sine[28408]=-66;
sine[28409]=-66;
sine[28410]=-66;
sine[28411]=-66;
sine[28412]=-66;
sine[28413]=-66;
sine[28414]=-66;
sine[28415]=-66;
sine[28416]=-66;
sine[28417]=-66;
sine[28418]=-65;
sine[28419]=-65;
sine[28420]=-65;
sine[28421]=-65;
sine[28422]=-65;
sine[28423]=-65;
sine[28424]=-65;
sine[28425]=-65;
sine[28426]=-65;
sine[28427]=-65;
sine[28428]=-65;
sine[28429]=-65;
sine[28430]=-65;
sine[28431]=-65;
sine[28432]=-65;
sine[28433]=-65;
sine[28434]=-65;
sine[28435]=-65;
sine[28436]=-65;
sine[28437]=-65;
sine[28438]=-65;
sine[28439]=-65;
sine[28440]=-65;
sine[28441]=-65;
sine[28442]=-65;
sine[28443]=-65;
sine[28444]=-65;
sine[28445]=-65;
sine[28446]=-65;
sine[28447]=-65;
sine[28448]=-65;
sine[28449]=-65;
sine[28450]=-65;
sine[28451]=-65;
sine[28452]=-65;
sine[28453]=-65;
sine[28454]=-65;
sine[28455]=-64;
sine[28456]=-64;
sine[28457]=-64;
sine[28458]=-64;
sine[28459]=-64;
sine[28460]=-64;
sine[28461]=-64;
sine[28462]=-64;
sine[28463]=-64;
sine[28464]=-64;
sine[28465]=-64;
sine[28466]=-64;
sine[28467]=-64;
sine[28468]=-64;
sine[28469]=-64;
sine[28470]=-64;
sine[28471]=-64;
sine[28472]=-64;
sine[28473]=-64;
sine[28474]=-64;
sine[28475]=-64;
sine[28476]=-64;
sine[28477]=-64;
sine[28478]=-64;
sine[28479]=-64;
sine[28480]=-64;
sine[28481]=-64;
sine[28482]=-64;
sine[28483]=-64;
sine[28484]=-64;
sine[28485]=-64;
sine[28486]=-64;
sine[28487]=-64;
sine[28488]=-64;
sine[28489]=-64;
sine[28490]=-63;
sine[28491]=-63;
sine[28492]=-63;
sine[28493]=-63;
sine[28494]=-63;
sine[28495]=-63;
sine[28496]=-63;
sine[28497]=-63;
sine[28498]=-63;
sine[28499]=-63;
sine[28500]=-63;
sine[28501]=-63;
sine[28502]=-63;
sine[28503]=-63;
sine[28504]=-63;
sine[28505]=-63;
sine[28506]=-63;
sine[28507]=-63;
sine[28508]=-63;
sine[28509]=-63;
sine[28510]=-63;
sine[28511]=-63;
sine[28512]=-63;
sine[28513]=-63;
sine[28514]=-63;
sine[28515]=-63;
sine[28516]=-63;
sine[28517]=-63;
sine[28518]=-63;
sine[28519]=-63;
sine[28520]=-63;
sine[28521]=-63;
sine[28522]=-63;
sine[28523]=-63;
sine[28524]=-63;
sine[28525]=-62;
sine[28526]=-62;
sine[28527]=-62;
sine[28528]=-62;
sine[28529]=-62;
sine[28530]=-62;
sine[28531]=-62;
sine[28532]=-62;
sine[28533]=-62;
sine[28534]=-62;
sine[28535]=-62;
sine[28536]=-62;
sine[28537]=-62;
sine[28538]=-62;
sine[28539]=-62;
sine[28540]=-62;
sine[28541]=-62;
sine[28542]=-62;
sine[28543]=-62;
sine[28544]=-62;
sine[28545]=-62;
sine[28546]=-62;
sine[28547]=-62;
sine[28548]=-62;
sine[28549]=-62;
sine[28550]=-62;
sine[28551]=-62;
sine[28552]=-62;
sine[28553]=-62;
sine[28554]=-62;
sine[28555]=-62;
sine[28556]=-62;
sine[28557]=-62;
sine[28558]=-61;
sine[28559]=-61;
sine[28560]=-61;
sine[28561]=-61;
sine[28562]=-61;
sine[28563]=-61;
sine[28564]=-61;
sine[28565]=-61;
sine[28566]=-61;
sine[28567]=-61;
sine[28568]=-61;
sine[28569]=-61;
sine[28570]=-61;
sine[28571]=-61;
sine[28572]=-61;
sine[28573]=-61;
sine[28574]=-61;
sine[28575]=-61;
sine[28576]=-61;
sine[28577]=-61;
sine[28578]=-61;
sine[28579]=-61;
sine[28580]=-61;
sine[28581]=-61;
sine[28582]=-61;
sine[28583]=-61;
sine[28584]=-61;
sine[28585]=-61;
sine[28586]=-61;
sine[28587]=-61;
sine[28588]=-61;
sine[28589]=-61;
sine[28590]=-61;
sine[28591]=-60;
sine[28592]=-60;
sine[28593]=-60;
sine[28594]=-60;
sine[28595]=-60;
sine[28596]=-60;
sine[28597]=-60;
sine[28598]=-60;
sine[28599]=-60;
sine[28600]=-60;
sine[28601]=-60;
sine[28602]=-60;
sine[28603]=-60;
sine[28604]=-60;
sine[28605]=-60;
sine[28606]=-60;
sine[28607]=-60;
sine[28608]=-60;
sine[28609]=-60;
sine[28610]=-60;
sine[28611]=-60;
sine[28612]=-60;
sine[28613]=-60;
sine[28614]=-60;
sine[28615]=-60;
sine[28616]=-60;
sine[28617]=-60;
sine[28618]=-60;
sine[28619]=-60;
sine[28620]=-60;
sine[28621]=-60;
sine[28622]=-60;
sine[28623]=-59;
sine[28624]=-59;
sine[28625]=-59;
sine[28626]=-59;
sine[28627]=-59;
sine[28628]=-59;
sine[28629]=-59;
sine[28630]=-59;
sine[28631]=-59;
sine[28632]=-59;
sine[28633]=-59;
sine[28634]=-59;
sine[28635]=-59;
sine[28636]=-59;
sine[28637]=-59;
sine[28638]=-59;
sine[28639]=-59;
sine[28640]=-59;
sine[28641]=-59;
sine[28642]=-59;
sine[28643]=-59;
sine[28644]=-59;
sine[28645]=-59;
sine[28646]=-59;
sine[28647]=-59;
sine[28648]=-59;
sine[28649]=-59;
sine[28650]=-59;
sine[28651]=-59;
sine[28652]=-59;
sine[28653]=-59;
sine[28654]=-58;
sine[28655]=-58;
sine[28656]=-58;
sine[28657]=-58;
sine[28658]=-58;
sine[28659]=-58;
sine[28660]=-58;
sine[28661]=-58;
sine[28662]=-58;
sine[28663]=-58;
sine[28664]=-58;
sine[28665]=-58;
sine[28666]=-58;
sine[28667]=-58;
sine[28668]=-58;
sine[28669]=-58;
sine[28670]=-58;
sine[28671]=-58;
sine[28672]=-58;
sine[28673]=-58;
sine[28674]=-58;
sine[28675]=-58;
sine[28676]=-58;
sine[28677]=-58;
sine[28678]=-58;
sine[28679]=-58;
sine[28680]=-58;
sine[28681]=-58;
sine[28682]=-58;
sine[28683]=-58;
sine[28684]=-57;
sine[28685]=-57;
sine[28686]=-57;
sine[28687]=-57;
sine[28688]=-57;
sine[28689]=-57;
sine[28690]=-57;
sine[28691]=-57;
sine[28692]=-57;
sine[28693]=-57;
sine[28694]=-57;
sine[28695]=-57;
sine[28696]=-57;
sine[28697]=-57;
sine[28698]=-57;
sine[28699]=-57;
sine[28700]=-57;
sine[28701]=-57;
sine[28702]=-57;
sine[28703]=-57;
sine[28704]=-57;
sine[28705]=-57;
sine[28706]=-57;
sine[28707]=-57;
sine[28708]=-57;
sine[28709]=-57;
sine[28710]=-57;
sine[28711]=-57;
sine[28712]=-57;
sine[28713]=-57;
sine[28714]=-56;
sine[28715]=-56;
sine[28716]=-56;
sine[28717]=-56;
sine[28718]=-56;
sine[28719]=-56;
sine[28720]=-56;
sine[28721]=-56;
sine[28722]=-56;
sine[28723]=-56;
sine[28724]=-56;
sine[28725]=-56;
sine[28726]=-56;
sine[28727]=-56;
sine[28728]=-56;
sine[28729]=-56;
sine[28730]=-56;
sine[28731]=-56;
sine[28732]=-56;
sine[28733]=-56;
sine[28734]=-56;
sine[28735]=-56;
sine[28736]=-56;
sine[28737]=-56;
sine[28738]=-56;
sine[28739]=-56;
sine[28740]=-56;
sine[28741]=-56;
sine[28742]=-56;
sine[28743]=-55;
sine[28744]=-55;
sine[28745]=-55;
sine[28746]=-55;
sine[28747]=-55;
sine[28748]=-55;
sine[28749]=-55;
sine[28750]=-55;
sine[28751]=-55;
sine[28752]=-55;
sine[28753]=-55;
sine[28754]=-55;
sine[28755]=-55;
sine[28756]=-55;
sine[28757]=-55;
sine[28758]=-55;
sine[28759]=-55;
sine[28760]=-55;
sine[28761]=-55;
sine[28762]=-55;
sine[28763]=-55;
sine[28764]=-55;
sine[28765]=-55;
sine[28766]=-55;
sine[28767]=-55;
sine[28768]=-55;
sine[28769]=-55;
sine[28770]=-55;
sine[28771]=-55;
sine[28772]=-54;
sine[28773]=-54;
sine[28774]=-54;
sine[28775]=-54;
sine[28776]=-54;
sine[28777]=-54;
sine[28778]=-54;
sine[28779]=-54;
sine[28780]=-54;
sine[28781]=-54;
sine[28782]=-54;
sine[28783]=-54;
sine[28784]=-54;
sine[28785]=-54;
sine[28786]=-54;
sine[28787]=-54;
sine[28788]=-54;
sine[28789]=-54;
sine[28790]=-54;
sine[28791]=-54;
sine[28792]=-54;
sine[28793]=-54;
sine[28794]=-54;
sine[28795]=-54;
sine[28796]=-54;
sine[28797]=-54;
sine[28798]=-54;
sine[28799]=-54;
sine[28800]=-53;
sine[28801]=-53;
sine[28802]=-53;
sine[28803]=-53;
sine[28804]=-53;
sine[28805]=-53;
sine[28806]=-53;
sine[28807]=-53;
sine[28808]=-53;
sine[28809]=-53;
sine[28810]=-53;
sine[28811]=-53;
sine[28812]=-53;
sine[28813]=-53;
sine[28814]=-53;
sine[28815]=-53;
sine[28816]=-53;
sine[28817]=-53;
sine[28818]=-53;
sine[28819]=-53;
sine[28820]=-53;
sine[28821]=-53;
sine[28822]=-53;
sine[28823]=-53;
sine[28824]=-53;
sine[28825]=-53;
sine[28826]=-53;
sine[28827]=-53;
sine[28828]=-52;
sine[28829]=-52;
sine[28830]=-52;
sine[28831]=-52;
sine[28832]=-52;
sine[28833]=-52;
sine[28834]=-52;
sine[28835]=-52;
sine[28836]=-52;
sine[28837]=-52;
sine[28838]=-52;
sine[28839]=-52;
sine[28840]=-52;
sine[28841]=-52;
sine[28842]=-52;
sine[28843]=-52;
sine[28844]=-52;
sine[28845]=-52;
sine[28846]=-52;
sine[28847]=-52;
sine[28848]=-52;
sine[28849]=-52;
sine[28850]=-52;
sine[28851]=-52;
sine[28852]=-52;
sine[28853]=-52;
sine[28854]=-52;
sine[28855]=-51;
sine[28856]=-51;
sine[28857]=-51;
sine[28858]=-51;
sine[28859]=-51;
sine[28860]=-51;
sine[28861]=-51;
sine[28862]=-51;
sine[28863]=-51;
sine[28864]=-51;
sine[28865]=-51;
sine[28866]=-51;
sine[28867]=-51;
sine[28868]=-51;
sine[28869]=-51;
sine[28870]=-51;
sine[28871]=-51;
sine[28872]=-51;
sine[28873]=-51;
sine[28874]=-51;
sine[28875]=-51;
sine[28876]=-51;
sine[28877]=-51;
sine[28878]=-51;
sine[28879]=-51;
sine[28880]=-51;
sine[28881]=-51;
sine[28882]=-50;
sine[28883]=-50;
sine[28884]=-50;
sine[28885]=-50;
sine[28886]=-50;
sine[28887]=-50;
sine[28888]=-50;
sine[28889]=-50;
sine[28890]=-50;
sine[28891]=-50;
sine[28892]=-50;
sine[28893]=-50;
sine[28894]=-50;
sine[28895]=-50;
sine[28896]=-50;
sine[28897]=-50;
sine[28898]=-50;
sine[28899]=-50;
sine[28900]=-50;
sine[28901]=-50;
sine[28902]=-50;
sine[28903]=-50;
sine[28904]=-50;
sine[28905]=-50;
sine[28906]=-50;
sine[28907]=-50;
sine[28908]=-49;
sine[28909]=-49;
sine[28910]=-49;
sine[28911]=-49;
sine[28912]=-49;
sine[28913]=-49;
sine[28914]=-49;
sine[28915]=-49;
sine[28916]=-49;
sine[28917]=-49;
sine[28918]=-49;
sine[28919]=-49;
sine[28920]=-49;
sine[28921]=-49;
sine[28922]=-49;
sine[28923]=-49;
sine[28924]=-49;
sine[28925]=-49;
sine[28926]=-49;
sine[28927]=-49;
sine[28928]=-49;
sine[28929]=-49;
sine[28930]=-49;
sine[28931]=-49;
sine[28932]=-49;
sine[28933]=-49;
sine[28934]=-49;
sine[28935]=-48;
sine[28936]=-48;
sine[28937]=-48;
sine[28938]=-48;
sine[28939]=-48;
sine[28940]=-48;
sine[28941]=-48;
sine[28942]=-48;
sine[28943]=-48;
sine[28944]=-48;
sine[28945]=-48;
sine[28946]=-48;
sine[28947]=-48;
sine[28948]=-48;
sine[28949]=-48;
sine[28950]=-48;
sine[28951]=-48;
sine[28952]=-48;
sine[28953]=-48;
sine[28954]=-48;
sine[28955]=-48;
sine[28956]=-48;
sine[28957]=-48;
sine[28958]=-48;
sine[28959]=-48;
sine[28960]=-47;
sine[28961]=-47;
sine[28962]=-47;
sine[28963]=-47;
sine[28964]=-47;
sine[28965]=-47;
sine[28966]=-47;
sine[28967]=-47;
sine[28968]=-47;
sine[28969]=-47;
sine[28970]=-47;
sine[28971]=-47;
sine[28972]=-47;
sine[28973]=-47;
sine[28974]=-47;
sine[28975]=-47;
sine[28976]=-47;
sine[28977]=-47;
sine[28978]=-47;
sine[28979]=-47;
sine[28980]=-47;
sine[28981]=-47;
sine[28982]=-47;
sine[28983]=-47;
sine[28984]=-47;
sine[28985]=-47;
sine[28986]=-46;
sine[28987]=-46;
sine[28988]=-46;
sine[28989]=-46;
sine[28990]=-46;
sine[28991]=-46;
sine[28992]=-46;
sine[28993]=-46;
sine[28994]=-46;
sine[28995]=-46;
sine[28996]=-46;
sine[28997]=-46;
sine[28998]=-46;
sine[28999]=-46;
sine[29000]=-46;
sine[29001]=-46;
sine[29002]=-46;
sine[29003]=-46;
sine[29004]=-46;
sine[29005]=-46;
sine[29006]=-46;
sine[29007]=-46;
sine[29008]=-46;
sine[29009]=-46;
sine[29010]=-46;
sine[29011]=-45;
sine[29012]=-45;
sine[29013]=-45;
sine[29014]=-45;
sine[29015]=-45;
sine[29016]=-45;
sine[29017]=-45;
sine[29018]=-45;
sine[29019]=-45;
sine[29020]=-45;
sine[29021]=-45;
sine[29022]=-45;
sine[29023]=-45;
sine[29024]=-45;
sine[29025]=-45;
sine[29026]=-45;
sine[29027]=-45;
sine[29028]=-45;
sine[29029]=-45;
sine[29030]=-45;
sine[29031]=-45;
sine[29032]=-45;
sine[29033]=-45;
sine[29034]=-45;
sine[29035]=-45;
sine[29036]=-44;
sine[29037]=-44;
sine[29038]=-44;
sine[29039]=-44;
sine[29040]=-44;
sine[29041]=-44;
sine[29042]=-44;
sine[29043]=-44;
sine[29044]=-44;
sine[29045]=-44;
sine[29046]=-44;
sine[29047]=-44;
sine[29048]=-44;
sine[29049]=-44;
sine[29050]=-44;
sine[29051]=-44;
sine[29052]=-44;
sine[29053]=-44;
sine[29054]=-44;
sine[29055]=-44;
sine[29056]=-44;
sine[29057]=-44;
sine[29058]=-44;
sine[29059]=-44;
sine[29060]=-44;
sine[29061]=-43;
sine[29062]=-43;
sine[29063]=-43;
sine[29064]=-43;
sine[29065]=-43;
sine[29066]=-43;
sine[29067]=-43;
sine[29068]=-43;
sine[29069]=-43;
sine[29070]=-43;
sine[29071]=-43;
sine[29072]=-43;
sine[29073]=-43;
sine[29074]=-43;
sine[29075]=-43;
sine[29076]=-43;
sine[29077]=-43;
sine[29078]=-43;
sine[29079]=-43;
sine[29080]=-43;
sine[29081]=-43;
sine[29082]=-43;
sine[29083]=-43;
sine[29084]=-43;
sine[29085]=-42;
sine[29086]=-42;
sine[29087]=-42;
sine[29088]=-42;
sine[29089]=-42;
sine[29090]=-42;
sine[29091]=-42;
sine[29092]=-42;
sine[29093]=-42;
sine[29094]=-42;
sine[29095]=-42;
sine[29096]=-42;
sine[29097]=-42;
sine[29098]=-42;
sine[29099]=-42;
sine[29100]=-42;
sine[29101]=-42;
sine[29102]=-42;
sine[29103]=-42;
sine[29104]=-42;
sine[29105]=-42;
sine[29106]=-42;
sine[29107]=-42;
sine[29108]=-42;
sine[29109]=-41;
sine[29110]=-41;
sine[29111]=-41;
sine[29112]=-41;
sine[29113]=-41;
sine[29114]=-41;
sine[29115]=-41;
sine[29116]=-41;
sine[29117]=-41;
sine[29118]=-41;
sine[29119]=-41;
sine[29120]=-41;
sine[29121]=-41;
sine[29122]=-41;
sine[29123]=-41;
sine[29124]=-41;
sine[29125]=-41;
sine[29126]=-41;
sine[29127]=-41;
sine[29128]=-41;
sine[29129]=-41;
sine[29130]=-41;
sine[29131]=-41;
sine[29132]=-41;
sine[29133]=-40;
sine[29134]=-40;
sine[29135]=-40;
sine[29136]=-40;
sine[29137]=-40;
sine[29138]=-40;
sine[29139]=-40;
sine[29140]=-40;
sine[29141]=-40;
sine[29142]=-40;
sine[29143]=-40;
sine[29144]=-40;
sine[29145]=-40;
sine[29146]=-40;
sine[29147]=-40;
sine[29148]=-40;
sine[29149]=-40;
sine[29150]=-40;
sine[29151]=-40;
sine[29152]=-40;
sine[29153]=-40;
sine[29154]=-40;
sine[29155]=-40;
sine[29156]=-40;
sine[29157]=-39;
sine[29158]=-39;
sine[29159]=-39;
sine[29160]=-39;
sine[29161]=-39;
sine[29162]=-39;
sine[29163]=-39;
sine[29164]=-39;
sine[29165]=-39;
sine[29166]=-39;
sine[29167]=-39;
sine[29168]=-39;
sine[29169]=-39;
sine[29170]=-39;
sine[29171]=-39;
sine[29172]=-39;
sine[29173]=-39;
sine[29174]=-39;
sine[29175]=-39;
sine[29176]=-39;
sine[29177]=-39;
sine[29178]=-39;
sine[29179]=-39;
sine[29180]=-38;
sine[29181]=-38;
sine[29182]=-38;
sine[29183]=-38;
sine[29184]=-38;
sine[29185]=-38;
sine[29186]=-38;
sine[29187]=-38;
sine[29188]=-38;
sine[29189]=-38;
sine[29190]=-38;
sine[29191]=-38;
sine[29192]=-38;
sine[29193]=-38;
sine[29194]=-38;
sine[29195]=-38;
sine[29196]=-38;
sine[29197]=-38;
sine[29198]=-38;
sine[29199]=-38;
sine[29200]=-38;
sine[29201]=-38;
sine[29202]=-38;
sine[29203]=-38;
sine[29204]=-37;
sine[29205]=-37;
sine[29206]=-37;
sine[29207]=-37;
sine[29208]=-37;
sine[29209]=-37;
sine[29210]=-37;
sine[29211]=-37;
sine[29212]=-37;
sine[29213]=-37;
sine[29214]=-37;
sine[29215]=-37;
sine[29216]=-37;
sine[29217]=-37;
sine[29218]=-37;
sine[29219]=-37;
sine[29220]=-37;
sine[29221]=-37;
sine[29222]=-37;
sine[29223]=-37;
sine[29224]=-37;
sine[29225]=-37;
sine[29226]=-37;
sine[29227]=-36;
sine[29228]=-36;
sine[29229]=-36;
sine[29230]=-36;
sine[29231]=-36;
sine[29232]=-36;
sine[29233]=-36;
sine[29234]=-36;
sine[29235]=-36;
sine[29236]=-36;
sine[29237]=-36;
sine[29238]=-36;
sine[29239]=-36;
sine[29240]=-36;
sine[29241]=-36;
sine[29242]=-36;
sine[29243]=-36;
sine[29244]=-36;
sine[29245]=-36;
sine[29246]=-36;
sine[29247]=-36;
sine[29248]=-36;
sine[29249]=-36;
sine[29250]=-35;
sine[29251]=-35;
sine[29252]=-35;
sine[29253]=-35;
sine[29254]=-35;
sine[29255]=-35;
sine[29256]=-35;
sine[29257]=-35;
sine[29258]=-35;
sine[29259]=-35;
sine[29260]=-35;
sine[29261]=-35;
sine[29262]=-35;
sine[29263]=-35;
sine[29264]=-35;
sine[29265]=-35;
sine[29266]=-35;
sine[29267]=-35;
sine[29268]=-35;
sine[29269]=-35;
sine[29270]=-35;
sine[29271]=-35;
sine[29272]=-35;
sine[29273]=-34;
sine[29274]=-34;
sine[29275]=-34;
sine[29276]=-34;
sine[29277]=-34;
sine[29278]=-34;
sine[29279]=-34;
sine[29280]=-34;
sine[29281]=-34;
sine[29282]=-34;
sine[29283]=-34;
sine[29284]=-34;
sine[29285]=-34;
sine[29286]=-34;
sine[29287]=-34;
sine[29288]=-34;
sine[29289]=-34;
sine[29290]=-34;
sine[29291]=-34;
sine[29292]=-34;
sine[29293]=-34;
sine[29294]=-34;
sine[29295]=-33;
sine[29296]=-33;
sine[29297]=-33;
sine[29298]=-33;
sine[29299]=-33;
sine[29300]=-33;
sine[29301]=-33;
sine[29302]=-33;
sine[29303]=-33;
sine[29304]=-33;
sine[29305]=-33;
sine[29306]=-33;
sine[29307]=-33;
sine[29308]=-33;
sine[29309]=-33;
sine[29310]=-33;
sine[29311]=-33;
sine[29312]=-33;
sine[29313]=-33;
sine[29314]=-33;
sine[29315]=-33;
sine[29316]=-33;
sine[29317]=-33;
sine[29318]=-32;
sine[29319]=-32;
sine[29320]=-32;
sine[29321]=-32;
sine[29322]=-32;
sine[29323]=-32;
sine[29324]=-32;
sine[29325]=-32;
sine[29326]=-32;
sine[29327]=-32;
sine[29328]=-32;
sine[29329]=-32;
sine[29330]=-32;
sine[29331]=-32;
sine[29332]=-32;
sine[29333]=-32;
sine[29334]=-32;
sine[29335]=-32;
sine[29336]=-32;
sine[29337]=-32;
sine[29338]=-32;
sine[29339]=-32;
sine[29340]=-31;
sine[29341]=-31;
sine[29342]=-31;
sine[29343]=-31;
sine[29344]=-31;
sine[29345]=-31;
sine[29346]=-31;
sine[29347]=-31;
sine[29348]=-31;
sine[29349]=-31;
sine[29350]=-31;
sine[29351]=-31;
sine[29352]=-31;
sine[29353]=-31;
sine[29354]=-31;
sine[29355]=-31;
sine[29356]=-31;
sine[29357]=-31;
sine[29358]=-31;
sine[29359]=-31;
sine[29360]=-31;
sine[29361]=-31;
sine[29362]=-30;
sine[29363]=-30;
sine[29364]=-30;
sine[29365]=-30;
sine[29366]=-30;
sine[29367]=-30;
sine[29368]=-30;
sine[29369]=-30;
sine[29370]=-30;
sine[29371]=-30;
sine[29372]=-30;
sine[29373]=-30;
sine[29374]=-30;
sine[29375]=-30;
sine[29376]=-30;
sine[29377]=-30;
sine[29378]=-30;
sine[29379]=-30;
sine[29380]=-30;
sine[29381]=-30;
sine[29382]=-30;
sine[29383]=-30;
sine[29384]=-29;
sine[29385]=-29;
sine[29386]=-29;
sine[29387]=-29;
sine[29388]=-29;
sine[29389]=-29;
sine[29390]=-29;
sine[29391]=-29;
sine[29392]=-29;
sine[29393]=-29;
sine[29394]=-29;
sine[29395]=-29;
sine[29396]=-29;
sine[29397]=-29;
sine[29398]=-29;
sine[29399]=-29;
sine[29400]=-29;
sine[29401]=-29;
sine[29402]=-29;
sine[29403]=-29;
sine[29404]=-29;
sine[29405]=-29;
sine[29406]=-28;
sine[29407]=-28;
sine[29408]=-28;
sine[29409]=-28;
sine[29410]=-28;
sine[29411]=-28;
sine[29412]=-28;
sine[29413]=-28;
sine[29414]=-28;
sine[29415]=-28;
sine[29416]=-28;
sine[29417]=-28;
sine[29418]=-28;
sine[29419]=-28;
sine[29420]=-28;
sine[29421]=-28;
sine[29422]=-28;
sine[29423]=-28;
sine[29424]=-28;
sine[29425]=-28;
sine[29426]=-28;
sine[29427]=-28;
sine[29428]=-27;
sine[29429]=-27;
sine[29430]=-27;
sine[29431]=-27;
sine[29432]=-27;
sine[29433]=-27;
sine[29434]=-27;
sine[29435]=-27;
sine[29436]=-27;
sine[29437]=-27;
sine[29438]=-27;
sine[29439]=-27;
sine[29440]=-27;
sine[29441]=-27;
sine[29442]=-27;
sine[29443]=-27;
sine[29444]=-27;
sine[29445]=-27;
sine[29446]=-27;
sine[29447]=-27;
sine[29448]=-27;
sine[29449]=-27;
sine[29450]=-26;
sine[29451]=-26;
sine[29452]=-26;
sine[29453]=-26;
sine[29454]=-26;
sine[29455]=-26;
sine[29456]=-26;
sine[29457]=-26;
sine[29458]=-26;
sine[29459]=-26;
sine[29460]=-26;
sine[29461]=-26;
sine[29462]=-26;
sine[29463]=-26;
sine[29464]=-26;
sine[29465]=-26;
sine[29466]=-26;
sine[29467]=-26;
sine[29468]=-26;
sine[29469]=-26;
sine[29470]=-26;
sine[29471]=-25;
sine[29472]=-25;
sine[29473]=-25;
sine[29474]=-25;
sine[29475]=-25;
sine[29476]=-25;
sine[29477]=-25;
sine[29478]=-25;
sine[29479]=-25;
sine[29480]=-25;
sine[29481]=-25;
sine[29482]=-25;
sine[29483]=-25;
sine[29484]=-25;
sine[29485]=-25;
sine[29486]=-25;
sine[29487]=-25;
sine[29488]=-25;
sine[29489]=-25;
sine[29490]=-25;
sine[29491]=-25;
sine[29492]=-25;
sine[29493]=-24;
sine[29494]=-24;
sine[29495]=-24;
sine[29496]=-24;
sine[29497]=-24;
sine[29498]=-24;
sine[29499]=-24;
sine[29500]=-24;
sine[29501]=-24;
sine[29502]=-24;
sine[29503]=-24;
sine[29504]=-24;
sine[29505]=-24;
sine[29506]=-24;
sine[29507]=-24;
sine[29508]=-24;
sine[29509]=-24;
sine[29510]=-24;
sine[29511]=-24;
sine[29512]=-24;
sine[29513]=-24;
sine[29514]=-23;
sine[29515]=-23;
sine[29516]=-23;
sine[29517]=-23;
sine[29518]=-23;
sine[29519]=-23;
sine[29520]=-23;
sine[29521]=-23;
sine[29522]=-23;
sine[29523]=-23;
sine[29524]=-23;
sine[29525]=-23;
sine[29526]=-23;
sine[29527]=-23;
sine[29528]=-23;
sine[29529]=-23;
sine[29530]=-23;
sine[29531]=-23;
sine[29532]=-23;
sine[29533]=-23;
sine[29534]=-23;
sine[29535]=-23;
sine[29536]=-22;
sine[29537]=-22;
sine[29538]=-22;
sine[29539]=-22;
sine[29540]=-22;
sine[29541]=-22;
sine[29542]=-22;
sine[29543]=-22;
sine[29544]=-22;
sine[29545]=-22;
sine[29546]=-22;
sine[29547]=-22;
sine[29548]=-22;
sine[29549]=-22;
sine[29550]=-22;
sine[29551]=-22;
sine[29552]=-22;
sine[29553]=-22;
sine[29554]=-22;
sine[29555]=-22;
sine[29556]=-22;
sine[29557]=-21;
sine[29558]=-21;
sine[29559]=-21;
sine[29560]=-21;
sine[29561]=-21;
sine[29562]=-21;
sine[29563]=-21;
sine[29564]=-21;
sine[29565]=-21;
sine[29566]=-21;
sine[29567]=-21;
sine[29568]=-21;
sine[29569]=-21;
sine[29570]=-21;
sine[29571]=-21;
sine[29572]=-21;
sine[29573]=-21;
sine[29574]=-21;
sine[29575]=-21;
sine[29576]=-21;
sine[29577]=-21;
sine[29578]=-20;
sine[29579]=-20;
sine[29580]=-20;
sine[29581]=-20;
sine[29582]=-20;
sine[29583]=-20;
sine[29584]=-20;
sine[29585]=-20;
sine[29586]=-20;
sine[29587]=-20;
sine[29588]=-20;
sine[29589]=-20;
sine[29590]=-20;
sine[29591]=-20;
sine[29592]=-20;
sine[29593]=-20;
sine[29594]=-20;
sine[29595]=-20;
sine[29596]=-20;
sine[29597]=-20;
sine[29598]=-20;
sine[29599]=-19;
sine[29600]=-19;
sine[29601]=-19;
sine[29602]=-19;
sine[29603]=-19;
sine[29604]=-19;
sine[29605]=-19;
sine[29606]=-19;
sine[29607]=-19;
sine[29608]=-19;
sine[29609]=-19;
sine[29610]=-19;
sine[29611]=-19;
sine[29612]=-19;
sine[29613]=-19;
sine[29614]=-19;
sine[29615]=-19;
sine[29616]=-19;
sine[29617]=-19;
sine[29618]=-19;
sine[29619]=-19;
sine[29620]=-18;
sine[29621]=-18;
sine[29622]=-18;
sine[29623]=-18;
sine[29624]=-18;
sine[29625]=-18;
sine[29626]=-18;
sine[29627]=-18;
sine[29628]=-18;
sine[29629]=-18;
sine[29630]=-18;
sine[29631]=-18;
sine[29632]=-18;
sine[29633]=-18;
sine[29634]=-18;
sine[29635]=-18;
sine[29636]=-18;
sine[29637]=-18;
sine[29638]=-18;
sine[29639]=-18;
sine[29640]=-18;
sine[29641]=-17;
sine[29642]=-17;
sine[29643]=-17;
sine[29644]=-17;
sine[29645]=-17;
sine[29646]=-17;
sine[29647]=-17;
sine[29648]=-17;
sine[29649]=-17;
sine[29650]=-17;
sine[29651]=-17;
sine[29652]=-17;
sine[29653]=-17;
sine[29654]=-17;
sine[29655]=-17;
sine[29656]=-17;
sine[29657]=-17;
sine[29658]=-17;
sine[29659]=-17;
sine[29660]=-17;
sine[29661]=-17;
sine[29662]=-16;
sine[29663]=-16;
sine[29664]=-16;
sine[29665]=-16;
sine[29666]=-16;
sine[29667]=-16;
sine[29668]=-16;
sine[29669]=-16;
sine[29670]=-16;
sine[29671]=-16;
sine[29672]=-16;
sine[29673]=-16;
sine[29674]=-16;
sine[29675]=-16;
sine[29676]=-16;
sine[29677]=-16;
sine[29678]=-16;
sine[29679]=-16;
sine[29680]=-16;
sine[29681]=-16;
sine[29682]=-16;
sine[29683]=-15;
sine[29684]=-15;
sine[29685]=-15;
sine[29686]=-15;
sine[29687]=-15;
sine[29688]=-15;
sine[29689]=-15;
sine[29690]=-15;
sine[29691]=-15;
sine[29692]=-15;
sine[29693]=-15;
sine[29694]=-15;
sine[29695]=-15;
sine[29696]=-15;
sine[29697]=-15;
sine[29698]=-15;
sine[29699]=-15;
sine[29700]=-15;
sine[29701]=-15;
sine[29702]=-15;
sine[29703]=-14;
sine[29704]=-14;
sine[29705]=-14;
sine[29706]=-14;
sine[29707]=-14;
sine[29708]=-14;
sine[29709]=-14;
sine[29710]=-14;
sine[29711]=-14;
sine[29712]=-14;
sine[29713]=-14;
sine[29714]=-14;
sine[29715]=-14;
sine[29716]=-14;
sine[29717]=-14;
sine[29718]=-14;
sine[29719]=-14;
sine[29720]=-14;
sine[29721]=-14;
sine[29722]=-14;
sine[29723]=-14;
sine[29724]=-13;
sine[29725]=-13;
sine[29726]=-13;
sine[29727]=-13;
sine[29728]=-13;
sine[29729]=-13;
sine[29730]=-13;
sine[29731]=-13;
sine[29732]=-13;
sine[29733]=-13;
sine[29734]=-13;
sine[29735]=-13;
sine[29736]=-13;
sine[29737]=-13;
sine[29738]=-13;
sine[29739]=-13;
sine[29740]=-13;
sine[29741]=-13;
sine[29742]=-13;
sine[29743]=-13;
sine[29744]=-13;
sine[29745]=-12;
sine[29746]=-12;
sine[29747]=-12;
sine[29748]=-12;
sine[29749]=-12;
sine[29750]=-12;
sine[29751]=-12;
sine[29752]=-12;
sine[29753]=-12;
sine[29754]=-12;
sine[29755]=-12;
sine[29756]=-12;
sine[29757]=-12;
sine[29758]=-12;
sine[29759]=-12;
sine[29760]=-12;
sine[29761]=-12;
sine[29762]=-12;
sine[29763]=-12;
sine[29764]=-12;
sine[29765]=-11;
sine[29766]=-11;
sine[29767]=-11;
sine[29768]=-11;
sine[29769]=-11;
sine[29770]=-11;
sine[29771]=-11;
sine[29772]=-11;
sine[29773]=-11;
sine[29774]=-11;
sine[29775]=-11;
sine[29776]=-11;
sine[29777]=-11;
sine[29778]=-11;
sine[29779]=-11;
sine[29780]=-11;
sine[29781]=-11;
sine[29782]=-11;
sine[29783]=-11;
sine[29784]=-11;
sine[29785]=-11;
sine[29786]=-10;
sine[29787]=-10;
sine[29788]=-10;
sine[29789]=-10;
sine[29790]=-10;
sine[29791]=-10;
sine[29792]=-10;
sine[29793]=-10;
sine[29794]=-10;
sine[29795]=-10;
sine[29796]=-10;
sine[29797]=-10;
sine[29798]=-10;
sine[29799]=-10;
sine[29800]=-10;
sine[29801]=-10;
sine[29802]=-10;
sine[29803]=-10;
sine[29804]=-10;
sine[29805]=-10;
sine[29806]=-9;
sine[29807]=-9;
sine[29808]=-9;
sine[29809]=-9;
sine[29810]=-9;
sine[29811]=-9;
sine[29812]=-9;
sine[29813]=-9;
sine[29814]=-9;
sine[29815]=-9;
sine[29816]=-9;
sine[29817]=-9;
sine[29818]=-9;
sine[29819]=-9;
sine[29820]=-9;
sine[29821]=-9;
sine[29822]=-9;
sine[29823]=-9;
sine[29824]=-9;
sine[29825]=-9;
sine[29826]=-9;
sine[29827]=-8;
sine[29828]=-8;
sine[29829]=-8;
sine[29830]=-8;
sine[29831]=-8;
sine[29832]=-8;
sine[29833]=-8;
sine[29834]=-8;
sine[29835]=-8;
sine[29836]=-8;
sine[29837]=-8;
sine[29838]=-8;
sine[29839]=-8;
sine[29840]=-8;
sine[29841]=-8;
sine[29842]=-8;
sine[29843]=-8;
sine[29844]=-8;
sine[29845]=-8;
sine[29846]=-8;
sine[29847]=-7;
sine[29848]=-7;
sine[29849]=-7;
sine[29850]=-7;
sine[29851]=-7;
sine[29852]=-7;
sine[29853]=-7;
sine[29854]=-7;
sine[29855]=-7;
sine[29856]=-7;
sine[29857]=-7;
sine[29858]=-7;
sine[29859]=-7;
sine[29860]=-7;
sine[29861]=-7;
sine[29862]=-7;
sine[29863]=-7;
sine[29864]=-7;
sine[29865]=-7;
sine[29866]=-7;
sine[29867]=-7;
sine[29868]=-6;
sine[29869]=-6;
sine[29870]=-6;
sine[29871]=-6;
sine[29872]=-6;
sine[29873]=-6;
sine[29874]=-6;
sine[29875]=-6;
sine[29876]=-6;
sine[29877]=-6;
sine[29878]=-6;
sine[29879]=-6;
sine[29880]=-6;
sine[29881]=-6;
sine[29882]=-6;
sine[29883]=-6;
sine[29884]=-6;
sine[29885]=-6;
sine[29886]=-6;
sine[29887]=-6;
sine[29888]=-5;
sine[29889]=-5;
sine[29890]=-5;
sine[29891]=-5;
sine[29892]=-5;
sine[29893]=-5;
sine[29894]=-5;
sine[29895]=-5;
sine[29896]=-5;
sine[29897]=-5;
sine[29898]=-5;
sine[29899]=-5;
sine[29900]=-5;
sine[29901]=-5;
sine[29902]=-5;
sine[29903]=-5;
sine[29904]=-5;
sine[29905]=-5;
sine[29906]=-5;
sine[29907]=-5;
sine[29908]=-5;
sine[29909]=-4;
sine[29910]=-4;
sine[29911]=-4;
sine[29912]=-4;
sine[29913]=-4;
sine[29914]=-4;
sine[29915]=-4;
sine[29916]=-4;
sine[29917]=-4;
sine[29918]=-4;
sine[29919]=-4;
sine[29920]=-4;
sine[29921]=-4;
sine[29922]=-4;
sine[29923]=-4;
sine[29924]=-4;
sine[29925]=-4;
sine[29926]=-4;
sine[29927]=-4;
sine[29928]=-4;
sine[29929]=-3;
sine[29930]=-3;
sine[29931]=-3;
sine[29932]=-3;
sine[29933]=-3;
sine[29934]=-3;
sine[29935]=-3;
sine[29936]=-3;
sine[29937]=-3;
sine[29938]=-3;
sine[29939]=-3;
sine[29940]=-3;
sine[29941]=-3;
sine[29942]=-3;
sine[29943]=-3;
sine[29944]=-3;
sine[29945]=-3;
sine[29946]=-3;
sine[29947]=-3;
sine[29948]=-3;
sine[29949]=-3;
sine[29950]=-2;
sine[29951]=-2;
sine[29952]=-2;
sine[29953]=-2;
sine[29954]=-2;
sine[29955]=-2;
sine[29956]=-2;
sine[29957]=-2;
sine[29958]=-2;
sine[29959]=-2;
sine[29960]=-2;
sine[29961]=-2;
sine[29962]=-2;
sine[29963]=-2;
sine[29964]=-2;
sine[29965]=-2;
sine[29966]=-2;
sine[29967]=-2;
sine[29968]=-2;
sine[29969]=-2;
sine[29970]=-1;
sine[29971]=-1;
sine[29972]=-1;
sine[29973]=-1;
sine[29974]=-1;
sine[29975]=-1;
sine[29976]=-1;
sine[29977]=-1;
sine[29978]=-1;
sine[29979]=-1;
sine[29980]=-1;
sine[29981]=-1;
sine[29982]=-1;
sine[29983]=-1;
sine[29984]=-1;
sine[29985]=-1;
sine[29986]=-1;
sine[29987]=-1;
sine[29988]=-1;
sine[29989]=-1;
sine[29990]=0;
sine[29991]=0;
sine[29992]=0;
sine[29993]=0;
sine[29994]=0;
sine[29995]=0;
sine[29996]=0;
sine[29997]=0;
sine[29998]=0;
sine[29999]=0;
sine[30000]=0;
sine[30001]=0;
sine[30002]=0;
sine[30003]=0;
sine[30004]=0;
sine[30005]=0;
sine[30006]=0;
sine[30007]=0;
sine[30008]=0;
sine[30009]=0;
sine[30010]=0;
sine[30011]=1;
sine[30012]=1;
sine[30013]=1;
sine[30014]=1;
sine[30015]=1;
sine[30016]=1;
sine[30017]=1;
sine[30018]=1;
sine[30019]=1;
sine[30020]=1;
sine[30021]=1;
sine[30022]=1;
sine[30023]=1;
sine[30024]=1;
sine[30025]=1;
sine[30026]=1;
sine[30027]=1;
sine[30028]=1;
sine[30029]=1;
sine[30030]=1;
sine[30031]=2;
sine[30032]=2;
sine[30033]=2;
sine[30034]=2;
sine[30035]=2;
sine[30036]=2;
sine[30037]=2;
sine[30038]=2;
sine[30039]=2;
sine[30040]=2;
sine[30041]=2;
sine[30042]=2;
sine[30043]=2;
sine[30044]=2;
sine[30045]=2;
sine[30046]=2;
sine[30047]=2;
sine[30048]=2;
sine[30049]=2;
sine[30050]=2;
sine[30051]=3;
sine[30052]=3;
sine[30053]=3;
sine[30054]=3;
sine[30055]=3;
sine[30056]=3;
sine[30057]=3;
sine[30058]=3;
sine[30059]=3;
sine[30060]=3;
sine[30061]=3;
sine[30062]=3;
sine[30063]=3;
sine[30064]=3;
sine[30065]=3;
sine[30066]=3;
sine[30067]=3;
sine[30068]=3;
sine[30069]=3;
sine[30070]=3;
sine[30071]=3;
sine[30072]=4;
sine[30073]=4;
sine[30074]=4;
sine[30075]=4;
sine[30076]=4;
sine[30077]=4;
sine[30078]=4;
sine[30079]=4;
sine[30080]=4;
sine[30081]=4;
sine[30082]=4;
sine[30083]=4;
sine[30084]=4;
sine[30085]=4;
sine[30086]=4;
sine[30087]=4;
sine[30088]=4;
sine[30089]=4;
sine[30090]=4;
sine[30091]=4;
sine[30092]=5;
sine[30093]=5;
sine[30094]=5;
sine[30095]=5;
sine[30096]=5;
sine[30097]=5;
sine[30098]=5;
sine[30099]=5;
sine[30100]=5;
sine[30101]=5;
sine[30102]=5;
sine[30103]=5;
sine[30104]=5;
sine[30105]=5;
sine[30106]=5;
sine[30107]=5;
sine[30108]=5;
sine[30109]=5;
sine[30110]=5;
sine[30111]=5;
sine[30112]=5;
sine[30113]=6;
sine[30114]=6;
sine[30115]=6;
sine[30116]=6;
sine[30117]=6;
sine[30118]=6;
sine[30119]=6;
sine[30120]=6;
sine[30121]=6;
sine[30122]=6;
sine[30123]=6;
sine[30124]=6;
sine[30125]=6;
sine[30126]=6;
sine[30127]=6;
sine[30128]=6;
sine[30129]=6;
sine[30130]=6;
sine[30131]=6;
sine[30132]=6;
sine[30133]=7;
sine[30134]=7;
sine[30135]=7;
sine[30136]=7;
sine[30137]=7;
sine[30138]=7;
sine[30139]=7;
sine[30140]=7;
sine[30141]=7;
sine[30142]=7;
sine[30143]=7;
sine[30144]=7;
sine[30145]=7;
sine[30146]=7;
sine[30147]=7;
sine[30148]=7;
sine[30149]=7;
sine[30150]=7;
sine[30151]=7;
sine[30152]=7;
sine[30153]=7;
sine[30154]=8;
sine[30155]=8;
sine[30156]=8;
sine[30157]=8;
sine[30158]=8;
sine[30159]=8;
sine[30160]=8;
sine[30161]=8;
sine[30162]=8;
sine[30163]=8;
sine[30164]=8;
sine[30165]=8;
sine[30166]=8;
sine[30167]=8;
sine[30168]=8;
sine[30169]=8;
sine[30170]=8;
sine[30171]=8;
sine[30172]=8;
sine[30173]=8;
sine[30174]=9;
sine[30175]=9;
sine[30176]=9;
sine[30177]=9;
sine[30178]=9;
sine[30179]=9;
sine[30180]=9;
sine[30181]=9;
sine[30182]=9;
sine[30183]=9;
sine[30184]=9;
sine[30185]=9;
sine[30186]=9;
sine[30187]=9;
sine[30188]=9;
sine[30189]=9;
sine[30190]=9;
sine[30191]=9;
sine[30192]=9;
sine[30193]=9;
sine[30194]=9;
sine[30195]=10;
sine[30196]=10;
sine[30197]=10;
sine[30198]=10;
sine[30199]=10;
sine[30200]=10;
sine[30201]=10;
sine[30202]=10;
sine[30203]=10;
sine[30204]=10;
sine[30205]=10;
sine[30206]=10;
sine[30207]=10;
sine[30208]=10;
sine[30209]=10;
sine[30210]=10;
sine[30211]=10;
sine[30212]=10;
sine[30213]=10;
sine[30214]=10;
sine[30215]=11;
sine[30216]=11;
sine[30217]=11;
sine[30218]=11;
sine[30219]=11;
sine[30220]=11;
sine[30221]=11;
sine[30222]=11;
sine[30223]=11;
sine[30224]=11;
sine[30225]=11;
sine[30226]=11;
sine[30227]=11;
sine[30228]=11;
sine[30229]=11;
sine[30230]=11;
sine[30231]=11;
sine[30232]=11;
sine[30233]=11;
sine[30234]=11;
sine[30235]=11;
sine[30236]=12;
sine[30237]=12;
sine[30238]=12;
sine[30239]=12;
sine[30240]=12;
sine[30241]=12;
sine[30242]=12;
sine[30243]=12;
sine[30244]=12;
sine[30245]=12;
sine[30246]=12;
sine[30247]=12;
sine[30248]=12;
sine[30249]=12;
sine[30250]=12;
sine[30251]=12;
sine[30252]=12;
sine[30253]=12;
sine[30254]=12;
sine[30255]=12;
sine[30256]=13;
sine[30257]=13;
sine[30258]=13;
sine[30259]=13;
sine[30260]=13;
sine[30261]=13;
sine[30262]=13;
sine[30263]=13;
sine[30264]=13;
sine[30265]=13;
sine[30266]=13;
sine[30267]=13;
sine[30268]=13;
sine[30269]=13;
sine[30270]=13;
sine[30271]=13;
sine[30272]=13;
sine[30273]=13;
sine[30274]=13;
sine[30275]=13;
sine[30276]=13;
sine[30277]=14;
sine[30278]=14;
sine[30279]=14;
sine[30280]=14;
sine[30281]=14;
sine[30282]=14;
sine[30283]=14;
sine[30284]=14;
sine[30285]=14;
sine[30286]=14;
sine[30287]=14;
sine[30288]=14;
sine[30289]=14;
sine[30290]=14;
sine[30291]=14;
sine[30292]=14;
sine[30293]=14;
sine[30294]=14;
sine[30295]=14;
sine[30296]=14;
sine[30297]=14;
sine[30298]=15;
sine[30299]=15;
sine[30300]=15;
sine[30301]=15;
sine[30302]=15;
sine[30303]=15;
sine[30304]=15;
sine[30305]=15;
sine[30306]=15;
sine[30307]=15;
sine[30308]=15;
sine[30309]=15;
sine[30310]=15;
sine[30311]=15;
sine[30312]=15;
sine[30313]=15;
sine[30314]=15;
sine[30315]=15;
sine[30316]=15;
sine[30317]=15;
sine[30318]=16;
sine[30319]=16;
sine[30320]=16;
sine[30321]=16;
sine[30322]=16;
sine[30323]=16;
sine[30324]=16;
sine[30325]=16;
sine[30326]=16;
sine[30327]=16;
sine[30328]=16;
sine[30329]=16;
sine[30330]=16;
sine[30331]=16;
sine[30332]=16;
sine[30333]=16;
sine[30334]=16;
sine[30335]=16;
sine[30336]=16;
sine[30337]=16;
sine[30338]=16;
sine[30339]=17;
sine[30340]=17;
sine[30341]=17;
sine[30342]=17;
sine[30343]=17;
sine[30344]=17;
sine[30345]=17;
sine[30346]=17;
sine[30347]=17;
sine[30348]=17;
sine[30349]=17;
sine[30350]=17;
sine[30351]=17;
sine[30352]=17;
sine[30353]=17;
sine[30354]=17;
sine[30355]=17;
sine[30356]=17;
sine[30357]=17;
sine[30358]=17;
sine[30359]=17;
sine[30360]=18;
sine[30361]=18;
sine[30362]=18;
sine[30363]=18;
sine[30364]=18;
sine[30365]=18;
sine[30366]=18;
sine[30367]=18;
sine[30368]=18;
sine[30369]=18;
sine[30370]=18;
sine[30371]=18;
sine[30372]=18;
sine[30373]=18;
sine[30374]=18;
sine[30375]=18;
sine[30376]=18;
sine[30377]=18;
sine[30378]=18;
sine[30379]=18;
sine[30380]=18;
sine[30381]=19;
sine[30382]=19;
sine[30383]=19;
sine[30384]=19;
sine[30385]=19;
sine[30386]=19;
sine[30387]=19;
sine[30388]=19;
sine[30389]=19;
sine[30390]=19;
sine[30391]=19;
sine[30392]=19;
sine[30393]=19;
sine[30394]=19;
sine[30395]=19;
sine[30396]=19;
sine[30397]=19;
sine[30398]=19;
sine[30399]=19;
sine[30400]=19;
sine[30401]=19;
sine[30402]=20;
sine[30403]=20;
sine[30404]=20;
sine[30405]=20;
sine[30406]=20;
sine[30407]=20;
sine[30408]=20;
sine[30409]=20;
sine[30410]=20;
sine[30411]=20;
sine[30412]=20;
sine[30413]=20;
sine[30414]=20;
sine[30415]=20;
sine[30416]=20;
sine[30417]=20;
sine[30418]=20;
sine[30419]=20;
sine[30420]=20;
sine[30421]=20;
sine[30422]=20;
sine[30423]=21;
sine[30424]=21;
sine[30425]=21;
sine[30426]=21;
sine[30427]=21;
sine[30428]=21;
sine[30429]=21;
sine[30430]=21;
sine[30431]=21;
sine[30432]=21;
sine[30433]=21;
sine[30434]=21;
sine[30435]=21;
sine[30436]=21;
sine[30437]=21;
sine[30438]=21;
sine[30439]=21;
sine[30440]=21;
sine[30441]=21;
sine[30442]=21;
sine[30443]=21;
sine[30444]=22;
sine[30445]=22;
sine[30446]=22;
sine[30447]=22;
sine[30448]=22;
sine[30449]=22;
sine[30450]=22;
sine[30451]=22;
sine[30452]=22;
sine[30453]=22;
sine[30454]=22;
sine[30455]=22;
sine[30456]=22;
sine[30457]=22;
sine[30458]=22;
sine[30459]=22;
sine[30460]=22;
sine[30461]=22;
sine[30462]=22;
sine[30463]=22;
sine[30464]=22;
sine[30465]=23;
sine[30466]=23;
sine[30467]=23;
sine[30468]=23;
sine[30469]=23;
sine[30470]=23;
sine[30471]=23;
sine[30472]=23;
sine[30473]=23;
sine[30474]=23;
sine[30475]=23;
sine[30476]=23;
sine[30477]=23;
sine[30478]=23;
sine[30479]=23;
sine[30480]=23;
sine[30481]=23;
sine[30482]=23;
sine[30483]=23;
sine[30484]=23;
sine[30485]=23;
sine[30486]=23;
sine[30487]=24;
sine[30488]=24;
sine[30489]=24;
sine[30490]=24;
sine[30491]=24;
sine[30492]=24;
sine[30493]=24;
sine[30494]=24;
sine[30495]=24;
sine[30496]=24;
sine[30497]=24;
sine[30498]=24;
sine[30499]=24;
sine[30500]=24;
sine[30501]=24;
sine[30502]=24;
sine[30503]=24;
sine[30504]=24;
sine[30505]=24;
sine[30506]=24;
sine[30507]=24;
sine[30508]=25;
sine[30509]=25;
sine[30510]=25;
sine[30511]=25;
sine[30512]=25;
sine[30513]=25;
sine[30514]=25;
sine[30515]=25;
sine[30516]=25;
sine[30517]=25;
sine[30518]=25;
sine[30519]=25;
sine[30520]=25;
sine[30521]=25;
sine[30522]=25;
sine[30523]=25;
sine[30524]=25;
sine[30525]=25;
sine[30526]=25;
sine[30527]=25;
sine[30528]=25;
sine[30529]=25;
sine[30530]=26;
sine[30531]=26;
sine[30532]=26;
sine[30533]=26;
sine[30534]=26;
sine[30535]=26;
sine[30536]=26;
sine[30537]=26;
sine[30538]=26;
sine[30539]=26;
sine[30540]=26;
sine[30541]=26;
sine[30542]=26;
sine[30543]=26;
sine[30544]=26;
sine[30545]=26;
sine[30546]=26;
sine[30547]=26;
sine[30548]=26;
sine[30549]=26;
sine[30550]=26;
sine[30551]=27;
sine[30552]=27;
sine[30553]=27;
sine[30554]=27;
sine[30555]=27;
sine[30556]=27;
sine[30557]=27;
sine[30558]=27;
sine[30559]=27;
sine[30560]=27;
sine[30561]=27;
sine[30562]=27;
sine[30563]=27;
sine[30564]=27;
sine[30565]=27;
sine[30566]=27;
sine[30567]=27;
sine[30568]=27;
sine[30569]=27;
sine[30570]=27;
sine[30571]=27;
sine[30572]=27;
sine[30573]=28;
sine[30574]=28;
sine[30575]=28;
sine[30576]=28;
sine[30577]=28;
sine[30578]=28;
sine[30579]=28;
sine[30580]=28;
sine[30581]=28;
sine[30582]=28;
sine[30583]=28;
sine[30584]=28;
sine[30585]=28;
sine[30586]=28;
sine[30587]=28;
sine[30588]=28;
sine[30589]=28;
sine[30590]=28;
sine[30591]=28;
sine[30592]=28;
sine[30593]=28;
sine[30594]=28;
sine[30595]=29;
sine[30596]=29;
sine[30597]=29;
sine[30598]=29;
sine[30599]=29;
sine[30600]=29;
sine[30601]=29;
sine[30602]=29;
sine[30603]=29;
sine[30604]=29;
sine[30605]=29;
sine[30606]=29;
sine[30607]=29;
sine[30608]=29;
sine[30609]=29;
sine[30610]=29;
sine[30611]=29;
sine[30612]=29;
sine[30613]=29;
sine[30614]=29;
sine[30615]=29;
sine[30616]=29;
sine[30617]=30;
sine[30618]=30;
sine[30619]=30;
sine[30620]=30;
sine[30621]=30;
sine[30622]=30;
sine[30623]=30;
sine[30624]=30;
sine[30625]=30;
sine[30626]=30;
sine[30627]=30;
sine[30628]=30;
sine[30629]=30;
sine[30630]=30;
sine[30631]=30;
sine[30632]=30;
sine[30633]=30;
sine[30634]=30;
sine[30635]=30;
sine[30636]=30;
sine[30637]=30;
sine[30638]=30;
sine[30639]=31;
sine[30640]=31;
sine[30641]=31;
sine[30642]=31;
sine[30643]=31;
sine[30644]=31;
sine[30645]=31;
sine[30646]=31;
sine[30647]=31;
sine[30648]=31;
sine[30649]=31;
sine[30650]=31;
sine[30651]=31;
sine[30652]=31;
sine[30653]=31;
sine[30654]=31;
sine[30655]=31;
sine[30656]=31;
sine[30657]=31;
sine[30658]=31;
sine[30659]=31;
sine[30660]=31;
sine[30661]=32;
sine[30662]=32;
sine[30663]=32;
sine[30664]=32;
sine[30665]=32;
sine[30666]=32;
sine[30667]=32;
sine[30668]=32;
sine[30669]=32;
sine[30670]=32;
sine[30671]=32;
sine[30672]=32;
sine[30673]=32;
sine[30674]=32;
sine[30675]=32;
sine[30676]=32;
sine[30677]=32;
sine[30678]=32;
sine[30679]=32;
sine[30680]=32;
sine[30681]=32;
sine[30682]=32;
sine[30683]=33;
sine[30684]=33;
sine[30685]=33;
sine[30686]=33;
sine[30687]=33;
sine[30688]=33;
sine[30689]=33;
sine[30690]=33;
sine[30691]=33;
sine[30692]=33;
sine[30693]=33;
sine[30694]=33;
sine[30695]=33;
sine[30696]=33;
sine[30697]=33;
sine[30698]=33;
sine[30699]=33;
sine[30700]=33;
sine[30701]=33;
sine[30702]=33;
sine[30703]=33;
sine[30704]=33;
sine[30705]=33;
sine[30706]=34;
sine[30707]=34;
sine[30708]=34;
sine[30709]=34;
sine[30710]=34;
sine[30711]=34;
sine[30712]=34;
sine[30713]=34;
sine[30714]=34;
sine[30715]=34;
sine[30716]=34;
sine[30717]=34;
sine[30718]=34;
sine[30719]=34;
sine[30720]=34;
sine[30721]=34;
sine[30722]=34;
sine[30723]=34;
sine[30724]=34;
sine[30725]=34;
sine[30726]=34;
sine[30727]=34;
sine[30728]=35;
sine[30729]=35;
sine[30730]=35;
sine[30731]=35;
sine[30732]=35;
sine[30733]=35;
sine[30734]=35;
sine[30735]=35;
sine[30736]=35;
sine[30737]=35;
sine[30738]=35;
sine[30739]=35;
sine[30740]=35;
sine[30741]=35;
sine[30742]=35;
sine[30743]=35;
sine[30744]=35;
sine[30745]=35;
sine[30746]=35;
sine[30747]=35;
sine[30748]=35;
sine[30749]=35;
sine[30750]=35;
sine[30751]=36;
sine[30752]=36;
sine[30753]=36;
sine[30754]=36;
sine[30755]=36;
sine[30756]=36;
sine[30757]=36;
sine[30758]=36;
sine[30759]=36;
sine[30760]=36;
sine[30761]=36;
sine[30762]=36;
sine[30763]=36;
sine[30764]=36;
sine[30765]=36;
sine[30766]=36;
sine[30767]=36;
sine[30768]=36;
sine[30769]=36;
sine[30770]=36;
sine[30771]=36;
sine[30772]=36;
sine[30773]=36;
sine[30774]=37;
sine[30775]=37;
sine[30776]=37;
sine[30777]=37;
sine[30778]=37;
sine[30779]=37;
sine[30780]=37;
sine[30781]=37;
sine[30782]=37;
sine[30783]=37;
sine[30784]=37;
sine[30785]=37;
sine[30786]=37;
sine[30787]=37;
sine[30788]=37;
sine[30789]=37;
sine[30790]=37;
sine[30791]=37;
sine[30792]=37;
sine[30793]=37;
sine[30794]=37;
sine[30795]=37;
sine[30796]=37;
sine[30797]=38;
sine[30798]=38;
sine[30799]=38;
sine[30800]=38;
sine[30801]=38;
sine[30802]=38;
sine[30803]=38;
sine[30804]=38;
sine[30805]=38;
sine[30806]=38;
sine[30807]=38;
sine[30808]=38;
sine[30809]=38;
sine[30810]=38;
sine[30811]=38;
sine[30812]=38;
sine[30813]=38;
sine[30814]=38;
sine[30815]=38;
sine[30816]=38;
sine[30817]=38;
sine[30818]=38;
sine[30819]=38;
sine[30820]=38;
sine[30821]=39;
sine[30822]=39;
sine[30823]=39;
sine[30824]=39;
sine[30825]=39;
sine[30826]=39;
sine[30827]=39;
sine[30828]=39;
sine[30829]=39;
sine[30830]=39;
sine[30831]=39;
sine[30832]=39;
sine[30833]=39;
sine[30834]=39;
sine[30835]=39;
sine[30836]=39;
sine[30837]=39;
sine[30838]=39;
sine[30839]=39;
sine[30840]=39;
sine[30841]=39;
sine[30842]=39;
sine[30843]=39;
sine[30844]=40;
sine[30845]=40;
sine[30846]=40;
sine[30847]=40;
sine[30848]=40;
sine[30849]=40;
sine[30850]=40;
sine[30851]=40;
sine[30852]=40;
sine[30853]=40;
sine[30854]=40;
sine[30855]=40;
sine[30856]=40;
sine[30857]=40;
sine[30858]=40;
sine[30859]=40;
sine[30860]=40;
sine[30861]=40;
sine[30862]=40;
sine[30863]=40;
sine[30864]=40;
sine[30865]=40;
sine[30866]=40;
sine[30867]=40;
sine[30868]=41;
sine[30869]=41;
sine[30870]=41;
sine[30871]=41;
sine[30872]=41;
sine[30873]=41;
sine[30874]=41;
sine[30875]=41;
sine[30876]=41;
sine[30877]=41;
sine[30878]=41;
sine[30879]=41;
sine[30880]=41;
sine[30881]=41;
sine[30882]=41;
sine[30883]=41;
sine[30884]=41;
sine[30885]=41;
sine[30886]=41;
sine[30887]=41;
sine[30888]=41;
sine[30889]=41;
sine[30890]=41;
sine[30891]=41;
sine[30892]=42;
sine[30893]=42;
sine[30894]=42;
sine[30895]=42;
sine[30896]=42;
sine[30897]=42;
sine[30898]=42;
sine[30899]=42;
sine[30900]=42;
sine[30901]=42;
sine[30902]=42;
sine[30903]=42;
sine[30904]=42;
sine[30905]=42;
sine[30906]=42;
sine[30907]=42;
sine[30908]=42;
sine[30909]=42;
sine[30910]=42;
sine[30911]=42;
sine[30912]=42;
sine[30913]=42;
sine[30914]=42;
sine[30915]=42;
sine[30916]=43;
sine[30917]=43;
sine[30918]=43;
sine[30919]=43;
sine[30920]=43;
sine[30921]=43;
sine[30922]=43;
sine[30923]=43;
sine[30924]=43;
sine[30925]=43;
sine[30926]=43;
sine[30927]=43;
sine[30928]=43;
sine[30929]=43;
sine[30930]=43;
sine[30931]=43;
sine[30932]=43;
sine[30933]=43;
sine[30934]=43;
sine[30935]=43;
sine[30936]=43;
sine[30937]=43;
sine[30938]=43;
sine[30939]=43;
sine[30940]=44;
sine[30941]=44;
sine[30942]=44;
sine[30943]=44;
sine[30944]=44;
sine[30945]=44;
sine[30946]=44;
sine[30947]=44;
sine[30948]=44;
sine[30949]=44;
sine[30950]=44;
sine[30951]=44;
sine[30952]=44;
sine[30953]=44;
sine[30954]=44;
sine[30955]=44;
sine[30956]=44;
sine[30957]=44;
sine[30958]=44;
sine[30959]=44;
sine[30960]=44;
sine[30961]=44;
sine[30962]=44;
sine[30963]=44;
sine[30964]=44;
sine[30965]=45;
sine[30966]=45;
sine[30967]=45;
sine[30968]=45;
sine[30969]=45;
sine[30970]=45;
sine[30971]=45;
sine[30972]=45;
sine[30973]=45;
sine[30974]=45;
sine[30975]=45;
sine[30976]=45;
sine[30977]=45;
sine[30978]=45;
sine[30979]=45;
sine[30980]=45;
sine[30981]=45;
sine[30982]=45;
sine[30983]=45;
sine[30984]=45;
sine[30985]=45;
sine[30986]=45;
sine[30987]=45;
sine[30988]=45;
sine[30989]=45;
sine[30990]=46;
sine[30991]=46;
sine[30992]=46;
sine[30993]=46;
sine[30994]=46;
sine[30995]=46;
sine[30996]=46;
sine[30997]=46;
sine[30998]=46;
sine[30999]=46;
sine[31000]=46;
sine[31001]=46;
sine[31002]=46;
sine[31003]=46;
sine[31004]=46;
sine[31005]=46;
sine[31006]=46;
sine[31007]=46;
sine[31008]=46;
sine[31009]=46;
sine[31010]=46;
sine[31011]=46;
sine[31012]=46;
sine[31013]=46;
sine[31014]=46;
sine[31015]=47;
sine[31016]=47;
sine[31017]=47;
sine[31018]=47;
sine[31019]=47;
sine[31020]=47;
sine[31021]=47;
sine[31022]=47;
sine[31023]=47;
sine[31024]=47;
sine[31025]=47;
sine[31026]=47;
sine[31027]=47;
sine[31028]=47;
sine[31029]=47;
sine[31030]=47;
sine[31031]=47;
sine[31032]=47;
sine[31033]=47;
sine[31034]=47;
sine[31035]=47;
sine[31036]=47;
sine[31037]=47;
sine[31038]=47;
sine[31039]=47;
sine[31040]=47;
sine[31041]=48;
sine[31042]=48;
sine[31043]=48;
sine[31044]=48;
sine[31045]=48;
sine[31046]=48;
sine[31047]=48;
sine[31048]=48;
sine[31049]=48;
sine[31050]=48;
sine[31051]=48;
sine[31052]=48;
sine[31053]=48;
sine[31054]=48;
sine[31055]=48;
sine[31056]=48;
sine[31057]=48;
sine[31058]=48;
sine[31059]=48;
sine[31060]=48;
sine[31061]=48;
sine[31062]=48;
sine[31063]=48;
sine[31064]=48;
sine[31065]=48;
sine[31066]=49;
sine[31067]=49;
sine[31068]=49;
sine[31069]=49;
sine[31070]=49;
sine[31071]=49;
sine[31072]=49;
sine[31073]=49;
sine[31074]=49;
sine[31075]=49;
sine[31076]=49;
sine[31077]=49;
sine[31078]=49;
sine[31079]=49;
sine[31080]=49;
sine[31081]=49;
sine[31082]=49;
sine[31083]=49;
sine[31084]=49;
sine[31085]=49;
sine[31086]=49;
sine[31087]=49;
sine[31088]=49;
sine[31089]=49;
sine[31090]=49;
sine[31091]=49;
sine[31092]=49;
sine[31093]=50;
sine[31094]=50;
sine[31095]=50;
sine[31096]=50;
sine[31097]=50;
sine[31098]=50;
sine[31099]=50;
sine[31100]=50;
sine[31101]=50;
sine[31102]=50;
sine[31103]=50;
sine[31104]=50;
sine[31105]=50;
sine[31106]=50;
sine[31107]=50;
sine[31108]=50;
sine[31109]=50;
sine[31110]=50;
sine[31111]=50;
sine[31112]=50;
sine[31113]=50;
sine[31114]=50;
sine[31115]=50;
sine[31116]=50;
sine[31117]=50;
sine[31118]=50;
sine[31119]=51;
sine[31120]=51;
sine[31121]=51;
sine[31122]=51;
sine[31123]=51;
sine[31124]=51;
sine[31125]=51;
sine[31126]=51;
sine[31127]=51;
sine[31128]=51;
sine[31129]=51;
sine[31130]=51;
sine[31131]=51;
sine[31132]=51;
sine[31133]=51;
sine[31134]=51;
sine[31135]=51;
sine[31136]=51;
sine[31137]=51;
sine[31138]=51;
sine[31139]=51;
sine[31140]=51;
sine[31141]=51;
sine[31142]=51;
sine[31143]=51;
sine[31144]=51;
sine[31145]=51;
sine[31146]=52;
sine[31147]=52;
sine[31148]=52;
sine[31149]=52;
sine[31150]=52;
sine[31151]=52;
sine[31152]=52;
sine[31153]=52;
sine[31154]=52;
sine[31155]=52;
sine[31156]=52;
sine[31157]=52;
sine[31158]=52;
sine[31159]=52;
sine[31160]=52;
sine[31161]=52;
sine[31162]=52;
sine[31163]=52;
sine[31164]=52;
sine[31165]=52;
sine[31166]=52;
sine[31167]=52;
sine[31168]=52;
sine[31169]=52;
sine[31170]=52;
sine[31171]=52;
sine[31172]=52;
sine[31173]=53;
sine[31174]=53;
sine[31175]=53;
sine[31176]=53;
sine[31177]=53;
sine[31178]=53;
sine[31179]=53;
sine[31180]=53;
sine[31181]=53;
sine[31182]=53;
sine[31183]=53;
sine[31184]=53;
sine[31185]=53;
sine[31186]=53;
sine[31187]=53;
sine[31188]=53;
sine[31189]=53;
sine[31190]=53;
sine[31191]=53;
sine[31192]=53;
sine[31193]=53;
sine[31194]=53;
sine[31195]=53;
sine[31196]=53;
sine[31197]=53;
sine[31198]=53;
sine[31199]=53;
sine[31200]=53;
sine[31201]=54;
sine[31202]=54;
sine[31203]=54;
sine[31204]=54;
sine[31205]=54;
sine[31206]=54;
sine[31207]=54;
sine[31208]=54;
sine[31209]=54;
sine[31210]=54;
sine[31211]=54;
sine[31212]=54;
sine[31213]=54;
sine[31214]=54;
sine[31215]=54;
sine[31216]=54;
sine[31217]=54;
sine[31218]=54;
sine[31219]=54;
sine[31220]=54;
sine[31221]=54;
sine[31222]=54;
sine[31223]=54;
sine[31224]=54;
sine[31225]=54;
sine[31226]=54;
sine[31227]=54;
sine[31228]=54;
sine[31229]=55;
sine[31230]=55;
sine[31231]=55;
sine[31232]=55;
sine[31233]=55;
sine[31234]=55;
sine[31235]=55;
sine[31236]=55;
sine[31237]=55;
sine[31238]=55;
sine[31239]=55;
sine[31240]=55;
sine[31241]=55;
sine[31242]=55;
sine[31243]=55;
sine[31244]=55;
sine[31245]=55;
sine[31246]=55;
sine[31247]=55;
sine[31248]=55;
sine[31249]=55;
sine[31250]=55;
sine[31251]=55;
sine[31252]=55;
sine[31253]=55;
sine[31254]=55;
sine[31255]=55;
sine[31256]=55;
sine[31257]=55;
sine[31258]=56;
sine[31259]=56;
sine[31260]=56;
sine[31261]=56;
sine[31262]=56;
sine[31263]=56;
sine[31264]=56;
sine[31265]=56;
sine[31266]=56;
sine[31267]=56;
sine[31268]=56;
sine[31269]=56;
sine[31270]=56;
sine[31271]=56;
sine[31272]=56;
sine[31273]=56;
sine[31274]=56;
sine[31275]=56;
sine[31276]=56;
sine[31277]=56;
sine[31278]=56;
sine[31279]=56;
sine[31280]=56;
sine[31281]=56;
sine[31282]=56;
sine[31283]=56;
sine[31284]=56;
sine[31285]=56;
sine[31286]=56;
sine[31287]=57;
sine[31288]=57;
sine[31289]=57;
sine[31290]=57;
sine[31291]=57;
sine[31292]=57;
sine[31293]=57;
sine[31294]=57;
sine[31295]=57;
sine[31296]=57;
sine[31297]=57;
sine[31298]=57;
sine[31299]=57;
sine[31300]=57;
sine[31301]=57;
sine[31302]=57;
sine[31303]=57;
sine[31304]=57;
sine[31305]=57;
sine[31306]=57;
sine[31307]=57;
sine[31308]=57;
sine[31309]=57;
sine[31310]=57;
sine[31311]=57;
sine[31312]=57;
sine[31313]=57;
sine[31314]=57;
sine[31315]=57;
sine[31316]=57;
sine[31317]=58;
sine[31318]=58;
sine[31319]=58;
sine[31320]=58;
sine[31321]=58;
sine[31322]=58;
sine[31323]=58;
sine[31324]=58;
sine[31325]=58;
sine[31326]=58;
sine[31327]=58;
sine[31328]=58;
sine[31329]=58;
sine[31330]=58;
sine[31331]=58;
sine[31332]=58;
sine[31333]=58;
sine[31334]=58;
sine[31335]=58;
sine[31336]=58;
sine[31337]=58;
sine[31338]=58;
sine[31339]=58;
sine[31340]=58;
sine[31341]=58;
sine[31342]=58;
sine[31343]=58;
sine[31344]=58;
sine[31345]=58;
sine[31346]=58;
sine[31347]=59;
sine[31348]=59;
sine[31349]=59;
sine[31350]=59;
sine[31351]=59;
sine[31352]=59;
sine[31353]=59;
sine[31354]=59;
sine[31355]=59;
sine[31356]=59;
sine[31357]=59;
sine[31358]=59;
sine[31359]=59;
sine[31360]=59;
sine[31361]=59;
sine[31362]=59;
sine[31363]=59;
sine[31364]=59;
sine[31365]=59;
sine[31366]=59;
sine[31367]=59;
sine[31368]=59;
sine[31369]=59;
sine[31370]=59;
sine[31371]=59;
sine[31372]=59;
sine[31373]=59;
sine[31374]=59;
sine[31375]=59;
sine[31376]=59;
sine[31377]=59;
sine[31378]=60;
sine[31379]=60;
sine[31380]=60;
sine[31381]=60;
sine[31382]=60;
sine[31383]=60;
sine[31384]=60;
sine[31385]=60;
sine[31386]=60;
sine[31387]=60;
sine[31388]=60;
sine[31389]=60;
sine[31390]=60;
sine[31391]=60;
sine[31392]=60;
sine[31393]=60;
sine[31394]=60;
sine[31395]=60;
sine[31396]=60;
sine[31397]=60;
sine[31398]=60;
sine[31399]=60;
sine[31400]=60;
sine[31401]=60;
sine[31402]=60;
sine[31403]=60;
sine[31404]=60;
sine[31405]=60;
sine[31406]=60;
sine[31407]=60;
sine[31408]=60;
sine[31409]=60;
sine[31410]=61;
sine[31411]=61;
sine[31412]=61;
sine[31413]=61;
sine[31414]=61;
sine[31415]=61;
sine[31416]=61;
sine[31417]=61;
sine[31418]=61;
sine[31419]=61;
sine[31420]=61;
sine[31421]=61;
sine[31422]=61;
sine[31423]=61;
sine[31424]=61;
sine[31425]=61;
sine[31426]=61;
sine[31427]=61;
sine[31428]=61;
sine[31429]=61;
sine[31430]=61;
sine[31431]=61;
sine[31432]=61;
sine[31433]=61;
sine[31434]=61;
sine[31435]=61;
sine[31436]=61;
sine[31437]=61;
sine[31438]=61;
sine[31439]=61;
sine[31440]=61;
sine[31441]=61;
sine[31442]=61;
sine[31443]=62;
sine[31444]=62;
sine[31445]=62;
sine[31446]=62;
sine[31447]=62;
sine[31448]=62;
sine[31449]=62;
sine[31450]=62;
sine[31451]=62;
sine[31452]=62;
sine[31453]=62;
sine[31454]=62;
sine[31455]=62;
sine[31456]=62;
sine[31457]=62;
sine[31458]=62;
sine[31459]=62;
sine[31460]=62;
sine[31461]=62;
sine[31462]=62;
sine[31463]=62;
sine[31464]=62;
sine[31465]=62;
sine[31466]=62;
sine[31467]=62;
sine[31468]=62;
sine[31469]=62;
sine[31470]=62;
sine[31471]=62;
sine[31472]=62;
sine[31473]=62;
sine[31474]=62;
sine[31475]=62;
sine[31476]=63;
sine[31477]=63;
sine[31478]=63;
sine[31479]=63;
sine[31480]=63;
sine[31481]=63;
sine[31482]=63;
sine[31483]=63;
sine[31484]=63;
sine[31485]=63;
sine[31486]=63;
sine[31487]=63;
sine[31488]=63;
sine[31489]=63;
sine[31490]=63;
sine[31491]=63;
sine[31492]=63;
sine[31493]=63;
sine[31494]=63;
sine[31495]=63;
sine[31496]=63;
sine[31497]=63;
sine[31498]=63;
sine[31499]=63;
sine[31500]=63;
sine[31501]=63;
sine[31502]=63;
sine[31503]=63;
sine[31504]=63;
sine[31505]=63;
sine[31506]=63;
sine[31507]=63;
sine[31508]=63;
sine[31509]=63;
sine[31510]=63;
sine[31511]=64;
sine[31512]=64;
sine[31513]=64;
sine[31514]=64;
sine[31515]=64;
sine[31516]=64;
sine[31517]=64;
sine[31518]=64;
sine[31519]=64;
sine[31520]=64;
sine[31521]=64;
sine[31522]=64;
sine[31523]=64;
sine[31524]=64;
sine[31525]=64;
sine[31526]=64;
sine[31527]=64;
sine[31528]=64;
sine[31529]=64;
sine[31530]=64;
sine[31531]=64;
sine[31532]=64;
sine[31533]=64;
sine[31534]=64;
sine[31535]=64;
sine[31536]=64;
sine[31537]=64;
sine[31538]=64;
sine[31539]=64;
sine[31540]=64;
sine[31541]=64;
sine[31542]=64;
sine[31543]=64;
sine[31544]=64;
sine[31545]=64;
sine[31546]=65;
sine[31547]=65;
sine[31548]=65;
sine[31549]=65;
sine[31550]=65;
sine[31551]=65;
sine[31552]=65;
sine[31553]=65;
sine[31554]=65;
sine[31555]=65;
sine[31556]=65;
sine[31557]=65;
sine[31558]=65;
sine[31559]=65;
sine[31560]=65;
sine[31561]=65;
sine[31562]=65;
sine[31563]=65;
sine[31564]=65;
sine[31565]=65;
sine[31566]=65;
sine[31567]=65;
sine[31568]=65;
sine[31569]=65;
sine[31570]=65;
sine[31571]=65;
sine[31572]=65;
sine[31573]=65;
sine[31574]=65;
sine[31575]=65;
sine[31576]=65;
sine[31577]=65;
sine[31578]=65;
sine[31579]=65;
sine[31580]=65;
sine[31581]=65;
sine[31582]=65;
sine[31583]=66;
sine[31584]=66;
sine[31585]=66;
sine[31586]=66;
sine[31587]=66;
sine[31588]=66;
sine[31589]=66;
sine[31590]=66;
sine[31591]=66;
sine[31592]=66;
sine[31593]=66;
sine[31594]=66;
sine[31595]=66;
sine[31596]=66;
sine[31597]=66;
sine[31598]=66;
sine[31599]=66;
sine[31600]=66;
sine[31601]=66;
sine[31602]=66;
sine[31603]=66;
sine[31604]=66;
sine[31605]=66;
sine[31606]=66;
sine[31607]=66;
sine[31608]=66;
sine[31609]=66;
sine[31610]=66;
sine[31611]=66;
sine[31612]=66;
sine[31613]=66;
sine[31614]=66;
sine[31615]=66;
sine[31616]=66;
sine[31617]=66;
sine[31618]=66;
sine[31619]=66;
sine[31620]=66;
sine[31621]=67;
sine[31622]=67;
sine[31623]=67;
sine[31624]=67;
sine[31625]=67;
sine[31626]=67;
sine[31627]=67;
sine[31628]=67;
sine[31629]=67;
sine[31630]=67;
sine[31631]=67;
sine[31632]=67;
sine[31633]=67;
sine[31634]=67;
sine[31635]=67;
sine[31636]=67;
sine[31637]=67;
sine[31638]=67;
sine[31639]=67;
sine[31640]=67;
sine[31641]=67;
sine[31642]=67;
sine[31643]=67;
sine[31644]=67;
sine[31645]=67;
sine[31646]=67;
sine[31647]=67;
sine[31648]=67;
sine[31649]=67;
sine[31650]=67;
sine[31651]=67;
sine[31652]=67;
sine[31653]=67;
sine[31654]=67;
sine[31655]=67;
sine[31656]=67;
sine[31657]=67;
sine[31658]=67;
sine[31659]=67;
sine[31660]=67;
sine[31661]=68;
sine[31662]=68;
sine[31663]=68;
sine[31664]=68;
sine[31665]=68;
sine[31666]=68;
sine[31667]=68;
sine[31668]=68;
sine[31669]=68;
sine[31670]=68;
sine[31671]=68;
sine[31672]=68;
sine[31673]=68;
sine[31674]=68;
sine[31675]=68;
sine[31676]=68;
sine[31677]=68;
sine[31678]=68;
sine[31679]=68;
sine[31680]=68;
sine[31681]=68;
sine[31682]=68;
sine[31683]=68;
sine[31684]=68;
sine[31685]=68;
sine[31686]=68;
sine[31687]=68;
sine[31688]=68;
sine[31689]=68;
sine[31690]=68;
sine[31691]=68;
sine[31692]=68;
sine[31693]=68;
sine[31694]=68;
sine[31695]=68;
sine[31696]=68;
sine[31697]=68;
sine[31698]=68;
sine[31699]=68;
sine[31700]=68;
sine[31701]=68;
sine[31702]=69;
sine[31703]=69;
sine[31704]=69;
sine[31705]=69;
sine[31706]=69;
sine[31707]=69;
sine[31708]=69;
sine[31709]=69;
sine[31710]=69;
sine[31711]=69;
sine[31712]=69;
sine[31713]=69;
sine[31714]=69;
sine[31715]=69;
sine[31716]=69;
sine[31717]=69;
sine[31718]=69;
sine[31719]=69;
sine[31720]=69;
sine[31721]=69;
sine[31722]=69;
sine[31723]=69;
sine[31724]=69;
sine[31725]=69;
sine[31726]=69;
sine[31727]=69;
sine[31728]=69;
sine[31729]=69;
sine[31730]=69;
sine[31731]=69;
sine[31732]=69;
sine[31733]=69;
sine[31734]=69;
sine[31735]=69;
sine[31736]=69;
sine[31737]=69;
sine[31738]=69;
sine[31739]=69;
sine[31740]=69;
sine[31741]=69;
sine[31742]=69;
sine[31743]=69;
sine[31744]=69;
sine[31745]=69;
sine[31746]=70;
sine[31747]=70;
sine[31748]=70;
sine[31749]=70;
sine[31750]=70;
sine[31751]=70;
sine[31752]=70;
sine[31753]=70;
sine[31754]=70;
sine[31755]=70;
sine[31756]=70;
sine[31757]=70;
sine[31758]=70;
sine[31759]=70;
sine[31760]=70;
sine[31761]=70;
sine[31762]=70;
sine[31763]=70;
sine[31764]=70;
sine[31765]=70;
sine[31766]=70;
sine[31767]=70;
sine[31768]=70;
sine[31769]=70;
sine[31770]=70;
sine[31771]=70;
sine[31772]=70;
sine[31773]=70;
sine[31774]=70;
sine[31775]=70;
sine[31776]=70;
sine[31777]=70;
sine[31778]=70;
sine[31779]=70;
sine[31780]=70;
sine[31781]=70;
sine[31782]=70;
sine[31783]=70;
sine[31784]=70;
sine[31785]=70;
sine[31786]=70;
sine[31787]=70;
sine[31788]=70;
sine[31789]=70;
sine[31790]=70;
sine[31791]=71;
sine[31792]=71;
sine[31793]=71;
sine[31794]=71;
sine[31795]=71;
sine[31796]=71;
sine[31797]=71;
sine[31798]=71;
sine[31799]=71;
sine[31800]=71;
sine[31801]=71;
sine[31802]=71;
sine[31803]=71;
sine[31804]=71;
sine[31805]=71;
sine[31806]=71;
sine[31807]=71;
sine[31808]=71;
sine[31809]=71;
sine[31810]=71;
sine[31811]=71;
sine[31812]=71;
sine[31813]=71;
sine[31814]=71;
sine[31815]=71;
sine[31816]=71;
sine[31817]=71;
sine[31818]=71;
sine[31819]=71;
sine[31820]=71;
sine[31821]=71;
sine[31822]=71;
sine[31823]=71;
sine[31824]=71;
sine[31825]=71;
sine[31826]=71;
sine[31827]=71;
sine[31828]=71;
sine[31829]=71;
sine[31830]=71;
sine[31831]=71;
sine[31832]=71;
sine[31833]=71;
sine[31834]=71;
sine[31835]=71;
sine[31836]=71;
sine[31837]=71;
sine[31838]=71;
sine[31839]=71;
sine[31840]=72;
sine[31841]=72;
sine[31842]=72;
sine[31843]=72;
sine[31844]=72;
sine[31845]=72;
sine[31846]=72;
sine[31847]=72;
sine[31848]=72;
sine[31849]=72;
sine[31850]=72;
sine[31851]=72;
sine[31852]=72;
sine[31853]=72;
sine[31854]=72;
sine[31855]=72;
sine[31856]=72;
sine[31857]=72;
sine[31858]=72;
sine[31859]=72;
sine[31860]=72;
sine[31861]=72;
sine[31862]=72;
sine[31863]=72;
sine[31864]=72;
sine[31865]=72;
sine[31866]=72;
sine[31867]=72;
sine[31868]=72;
sine[31869]=72;
sine[31870]=72;
sine[31871]=72;
sine[31872]=72;
sine[31873]=72;
sine[31874]=72;
sine[31875]=72;
sine[31876]=72;
sine[31877]=72;
sine[31878]=72;
sine[31879]=72;
sine[31880]=72;
sine[31881]=72;
sine[31882]=72;
sine[31883]=72;
sine[31884]=72;
sine[31885]=72;
sine[31886]=72;
sine[31887]=72;
sine[31888]=72;
sine[31889]=72;
sine[31890]=72;
sine[31891]=72;
sine[31892]=72;
sine[31893]=73;
sine[31894]=73;
sine[31895]=73;
sine[31896]=73;
sine[31897]=73;
sine[31898]=73;
sine[31899]=73;
sine[31900]=73;
sine[31901]=73;
sine[31902]=73;
sine[31903]=73;
sine[31904]=73;
sine[31905]=73;
sine[31906]=73;
sine[31907]=73;
sine[31908]=73;
sine[31909]=73;
sine[31910]=73;
sine[31911]=73;
sine[31912]=73;
sine[31913]=73;
sine[31914]=73;
sine[31915]=73;
sine[31916]=73;
sine[31917]=73;
sine[31918]=73;
sine[31919]=73;
sine[31920]=73;
sine[31921]=73;
sine[31922]=73;
sine[31923]=73;
sine[31924]=73;
sine[31925]=73;
sine[31926]=73;
sine[31927]=73;
sine[31928]=73;
sine[31929]=73;
sine[31930]=73;
sine[31931]=73;
sine[31932]=73;
sine[31933]=73;
sine[31934]=73;
sine[31935]=73;
sine[31936]=73;
sine[31937]=73;
sine[31938]=73;
sine[31939]=73;
sine[31940]=73;
sine[31941]=73;
sine[31942]=73;
sine[31943]=73;
sine[31944]=73;
sine[31945]=73;
sine[31946]=73;
sine[31947]=73;
sine[31948]=73;
sine[31949]=73;
sine[31950]=74;
sine[31951]=74;
sine[31952]=74;
sine[31953]=74;
sine[31954]=74;
sine[31955]=74;
sine[31956]=74;
sine[31957]=74;
sine[31958]=74;
sine[31959]=74;
sine[31960]=74;
sine[31961]=74;
sine[31962]=74;
sine[31963]=74;
sine[31964]=74;
sine[31965]=74;
sine[31966]=74;
sine[31967]=74;
sine[31968]=74;
sine[31969]=74;
sine[31970]=74;
sine[31971]=74;
sine[31972]=74;
sine[31973]=74;
sine[31974]=74;
sine[31975]=74;
sine[31976]=74;
sine[31977]=74;
sine[31978]=74;
sine[31979]=74;
sine[31980]=74;
sine[31981]=74;
sine[31982]=74;
sine[31983]=74;
sine[31984]=74;
sine[31985]=74;
sine[31986]=74;
sine[31987]=74;
sine[31988]=74;
sine[31989]=74;
sine[31990]=74;
sine[31991]=74;
sine[31992]=74;
sine[31993]=74;
sine[31994]=74;
sine[31995]=74;
sine[31996]=74;
sine[31997]=74;
sine[31998]=74;
sine[31999]=74;
sine[32000]=74;
sine[32001]=74;
sine[32002]=74;
sine[32003]=74;
sine[32004]=74;
sine[32005]=74;
sine[32006]=74;
sine[32007]=74;
sine[32008]=74;
sine[32009]=74;
sine[32010]=74;
sine[32011]=74;
sine[32012]=74;
sine[32013]=74;
sine[32014]=75;
sine[32015]=75;
sine[32016]=75;
sine[32017]=75;
sine[32018]=75;
sine[32019]=75;
sine[32020]=75;
sine[32021]=75;
sine[32022]=75;
sine[32023]=75;
sine[32024]=75;
sine[32025]=75;
sine[32026]=75;
sine[32027]=75;
sine[32028]=75;
sine[32029]=75;
sine[32030]=75;
sine[32031]=75;
sine[32032]=75;
sine[32033]=75;
sine[32034]=75;
sine[32035]=75;
sine[32036]=75;
sine[32037]=75;
sine[32038]=75;
sine[32039]=75;
sine[32040]=75;
sine[32041]=75;
sine[32042]=75;
sine[32043]=75;
sine[32044]=75;
sine[32045]=75;
sine[32046]=75;
sine[32047]=75;
sine[32048]=75;
sine[32049]=75;
sine[32050]=75;
sine[32051]=75;
sine[32052]=75;
sine[32053]=75;
sine[32054]=75;
sine[32055]=75;
sine[32056]=75;
sine[32057]=75;
sine[32058]=75;
sine[32059]=75;
sine[32060]=75;
sine[32061]=75;
sine[32062]=75;
sine[32063]=75;
sine[32064]=75;
sine[32065]=75;
sine[32066]=75;
sine[32067]=75;
sine[32068]=75;
sine[32069]=75;
sine[32070]=75;
sine[32071]=75;
sine[32072]=75;
sine[32073]=75;
sine[32074]=75;
sine[32075]=75;
sine[32076]=75;
sine[32077]=75;
sine[32078]=75;
sine[32079]=75;
sine[32080]=75;
sine[32081]=75;
sine[32082]=75;
sine[32083]=75;
sine[32084]=75;
sine[32085]=75;
sine[32086]=75;
sine[32087]=76;
sine[32088]=76;
sine[32089]=76;
sine[32090]=76;
sine[32091]=76;
sine[32092]=76;
sine[32093]=76;
sine[32094]=76;
sine[32095]=76;
sine[32096]=76;
sine[32097]=76;
sine[32098]=76;
sine[32099]=76;
sine[32100]=76;
sine[32101]=76;
sine[32102]=76;
sine[32103]=76;
sine[32104]=76;
sine[32105]=76;
sine[32106]=76;
sine[32107]=76;
sine[32108]=76;
sine[32109]=76;
sine[32110]=76;
sine[32111]=76;
sine[32112]=76;
sine[32113]=76;
sine[32114]=76;
sine[32115]=76;
sine[32116]=76;
sine[32117]=76;
sine[32118]=76;
sine[32119]=76;
sine[32120]=76;
sine[32121]=76;
sine[32122]=76;
sine[32123]=76;
sine[32124]=76;
sine[32125]=76;
sine[32126]=76;
sine[32127]=76;
sine[32128]=76;
sine[32129]=76;
sine[32130]=76;
sine[32131]=76;
sine[32132]=76;
sine[32133]=76;
sine[32134]=76;
sine[32135]=76;
sine[32136]=76;
sine[32137]=76;
sine[32138]=76;
sine[32139]=76;
sine[32140]=76;
sine[32141]=76;
sine[32142]=76;
sine[32143]=76;
sine[32144]=76;
sine[32145]=76;
sine[32146]=76;
sine[32147]=76;
sine[32148]=76;
sine[32149]=76;
sine[32150]=76;
sine[32151]=76;
sine[32152]=76;
sine[32153]=76;
sine[32154]=76;
sine[32155]=76;
sine[32156]=76;
sine[32157]=76;
sine[32158]=76;
sine[32159]=76;
sine[32160]=76;
sine[32161]=76;
sine[32162]=76;
sine[32163]=76;
sine[32164]=76;
sine[32165]=76;
sine[32166]=76;
sine[32167]=76;
sine[32168]=76;
sine[32169]=76;
sine[32170]=76;
sine[32171]=76;
sine[32172]=76;
sine[32173]=76;
sine[32174]=76;
sine[32175]=77;
sine[32176]=77;
sine[32177]=77;
sine[32178]=77;
sine[32179]=77;
sine[32180]=77;
sine[32181]=77;
sine[32182]=77;
sine[32183]=77;
sine[32184]=77;
sine[32185]=77;
sine[32186]=77;
sine[32187]=77;
sine[32188]=77;
sine[32189]=77;
sine[32190]=77;
sine[32191]=77;
sine[32192]=77;
sine[32193]=77;
sine[32194]=77;
sine[32195]=77;
sine[32196]=77;
sine[32197]=77;
sine[32198]=77;
sine[32199]=77;
sine[32200]=77;
sine[32201]=77;
sine[32202]=77;
sine[32203]=77;
sine[32204]=77;
sine[32205]=77;
sine[32206]=77;
sine[32207]=77;
sine[32208]=77;
sine[32209]=77;
sine[32210]=77;
sine[32211]=77;
sine[32212]=77;
sine[32213]=77;
sine[32214]=77;
sine[32215]=77;
sine[32216]=77;
sine[32217]=77;
sine[32218]=77;
sine[32219]=77;
sine[32220]=77;
sine[32221]=77;
sine[32222]=77;
sine[32223]=77;
sine[32224]=77;
sine[32225]=77;
sine[32226]=77;
sine[32227]=77;
sine[32228]=77;
sine[32229]=77;
sine[32230]=77;
sine[32231]=77;
sine[32232]=77;
sine[32233]=77;
sine[32234]=77;
sine[32235]=77;
sine[32236]=77;
sine[32237]=77;
sine[32238]=77;
sine[32239]=77;
sine[32240]=77;
sine[32241]=77;
sine[32242]=77;
sine[32243]=77;
sine[32244]=77;
sine[32245]=77;
sine[32246]=77;
sine[32247]=77;
sine[32248]=77;
sine[32249]=77;
sine[32250]=77;
sine[32251]=77;
sine[32252]=77;
sine[32253]=77;
sine[32254]=77;
sine[32255]=77;
sine[32256]=77;
sine[32257]=77;
sine[32258]=77;
sine[32259]=77;
sine[32260]=77;
sine[32261]=77;
sine[32262]=77;
sine[32263]=77;
sine[32264]=77;
sine[32265]=77;
sine[32266]=77;
sine[32267]=77;
sine[32268]=77;
sine[32269]=77;
sine[32270]=77;
sine[32271]=77;
sine[32272]=77;
sine[32273]=77;
sine[32274]=77;
sine[32275]=77;
sine[32276]=77;
sine[32277]=77;
sine[32278]=77;
sine[32279]=77;
sine[32280]=77;
sine[32281]=77;
sine[32282]=77;
sine[32283]=77;
sine[32284]=77;
sine[32285]=77;
sine[32286]=77;
sine[32287]=77;
sine[32288]=77;
sine[32289]=77;
sine[32290]=77;
sine[32291]=77;
sine[32292]=77;
sine[32293]=77;
sine[32294]=77;
sine[32295]=77;
sine[32296]=77;
sine[32297]=77;
sine[32298]=77;
sine[32299]=78;
sine[32300]=78;
sine[32301]=78;
sine[32302]=78;
sine[32303]=78;
sine[32304]=78;
sine[32305]=78;
sine[32306]=78;
sine[32307]=78;
sine[32308]=78;
sine[32309]=78;
sine[32310]=78;
sine[32311]=78;
sine[32312]=78;
sine[32313]=78;
sine[32314]=78;
sine[32315]=78;
sine[32316]=78;
sine[32317]=78;
sine[32318]=78;
sine[32319]=78;
sine[32320]=78;
sine[32321]=78;
sine[32322]=78;
sine[32323]=78;
sine[32324]=78;
sine[32325]=78;
sine[32326]=78;
sine[32327]=78;
sine[32328]=78;
sine[32329]=78;
sine[32330]=78;
sine[32331]=78;
sine[32332]=78;
sine[32333]=78;
sine[32334]=78;
sine[32335]=78;
sine[32336]=78;
sine[32337]=78;
sine[32338]=78;
sine[32339]=78;
sine[32340]=78;
sine[32341]=78;
sine[32342]=78;
sine[32343]=78;
sine[32344]=78;
sine[32345]=78;
sine[32346]=78;
sine[32347]=78;
sine[32348]=78;
sine[32349]=78;
sine[32350]=78;
sine[32351]=78;
sine[32352]=78;
sine[32353]=78;
sine[32354]=78;
sine[32355]=78;
sine[32356]=78;
sine[32357]=78;
sine[32358]=78;
sine[32359]=78;
sine[32360]=78;
sine[32361]=78;
sine[32362]=78;
sine[32363]=78;
sine[32364]=78;
sine[32365]=78;
sine[32366]=78;
sine[32367]=78;
sine[32368]=78;
sine[32369]=78;
sine[32370]=78;
sine[32371]=78;
sine[32372]=78;
sine[32373]=78;
sine[32374]=78;
sine[32375]=78;
sine[32376]=78;
sine[32377]=78;
sine[32378]=78;
sine[32379]=78;
sine[32380]=78;
sine[32381]=78;
sine[32382]=78;
sine[32383]=78;
sine[32384]=78;
sine[32385]=78;
sine[32386]=78;
sine[32387]=78;
sine[32388]=78;
sine[32389]=78;
sine[32390]=78;
sine[32391]=78;
sine[32392]=78;
sine[32393]=78;
sine[32394]=78;
sine[32395]=78;
sine[32396]=78;
sine[32397]=78;
sine[32398]=78;
sine[32399]=78;
sine[32400]=78;
sine[32401]=78;
sine[32402]=78;
sine[32403]=78;
sine[32404]=78;
sine[32405]=78;
sine[32406]=78;
sine[32407]=78;
sine[32408]=78;
sine[32409]=78;
sine[32410]=78;
sine[32411]=78;
sine[32412]=78;
sine[32413]=78;
sine[32414]=78;
sine[32415]=78;
sine[32416]=78;
sine[32417]=78;
sine[32418]=78;
sine[32419]=78;
sine[32420]=78;
sine[32421]=78;
sine[32422]=78;
sine[32423]=78;
sine[32424]=78;
sine[32425]=78;
sine[32426]=78;
sine[32427]=78;
sine[32428]=78;
sine[32429]=78;
sine[32430]=78;
sine[32431]=78;
sine[32432]=78;
sine[32433]=78;
sine[32434]=78;
sine[32435]=78;
sine[32436]=78;
sine[32437]=78;
sine[32438]=78;
sine[32439]=78;
sine[32440]=78;
sine[32441]=78;
sine[32442]=78;
sine[32443]=78;
sine[32444]=78;
sine[32445]=78;
sine[32446]=78;
sine[32447]=78;
sine[32448]=78;
sine[32449]=78;
sine[32450]=78;
sine[32451]=78;
sine[32452]=78;
sine[32453]=78;
sine[32454]=78;
sine[32455]=78;
sine[32456]=78;
sine[32457]=78;
sine[32458]=78;
sine[32459]=78;
sine[32460]=78;
sine[32461]=78;
sine[32462]=78;
sine[32463]=78;
sine[32464]=78;
sine[32465]=78;
sine[32466]=78;
sine[32467]=78;
sine[32468]=78;
sine[32469]=78;
sine[32470]=78;
sine[32471]=78;
sine[32472]=78;
sine[32473]=78;
sine[32474]=78;
sine[32475]=78;
sine[32476]=78;
sine[32477]=78;
sine[32478]=78;
sine[32479]=78;
sine[32480]=78;
sine[32481]=78;
sine[32482]=78;
sine[32483]=78;
sine[32484]=78;
sine[32485]=78;
sine[32486]=78;
sine[32487]=78;
sine[32488]=78;
sine[32489]=78;
sine[32490]=78;
sine[32491]=78;
sine[32492]=78;
sine[32493]=78;
sine[32494]=78;
sine[32495]=78;
sine[32496]=78;
sine[32497]=78;
sine[32498]=78;
sine[32499]=78;
sine[32500]=78;
sine[32501]=78;
sine[32502]=78;
sine[32503]=78;
sine[32504]=78;
sine[32505]=78;
sine[32506]=78;
sine[32507]=78;
sine[32508]=78;
sine[32509]=78;
sine[32510]=78;
sine[32511]=78;
sine[32512]=78;
sine[32513]=78;
sine[32514]=78;
sine[32515]=78;
sine[32516]=78;
sine[32517]=78;
sine[32518]=78;
sine[32519]=78;
sine[32520]=78;
sine[32521]=78;
sine[32522]=78;
sine[32523]=78;
sine[32524]=78;
sine[32525]=78;
sine[32526]=78;
sine[32527]=78;
sine[32528]=78;
sine[32529]=78;
sine[32530]=78;
sine[32531]=78;
sine[32532]=78;
sine[32533]=78;
sine[32534]=78;
sine[32535]=78;
sine[32536]=78;
sine[32537]=78;
sine[32538]=78;
sine[32539]=78;
sine[32540]=78;
sine[32541]=78;
sine[32542]=78;
sine[32543]=78;
sine[32544]=78;
sine[32545]=78;
sine[32546]=78;
sine[32547]=78;
sine[32548]=78;
sine[32549]=78;
sine[32550]=78;
sine[32551]=78;
sine[32552]=78;
sine[32553]=78;
sine[32554]=78;
sine[32555]=78;
sine[32556]=78;
sine[32557]=78;
sine[32558]=78;
sine[32559]=78;
sine[32560]=78;
sine[32561]=78;
sine[32562]=78;
sine[32563]=78;
sine[32564]=78;
sine[32565]=78;
sine[32566]=78;
sine[32567]=78;
sine[32568]=78;
sine[32569]=78;
sine[32570]=78;
sine[32571]=78;
sine[32572]=78;
sine[32573]=78;
sine[32574]=78;
sine[32575]=78;
sine[32576]=78;
sine[32577]=78;
sine[32578]=78;
sine[32579]=78;
sine[32580]=78;
sine[32581]=78;
sine[32582]=78;
sine[32583]=78;
sine[32584]=78;
sine[32585]=78;
sine[32586]=78;
sine[32587]=78;
sine[32588]=78;
sine[32589]=78;
sine[32590]=78;
sine[32591]=78;
sine[32592]=78;
sine[32593]=78;
sine[32594]=78;
sine[32595]=78;
sine[32596]=78;
sine[32597]=78;
sine[32598]=78;
sine[32599]=78;
sine[32600]=78;
sine[32601]=78;
sine[32602]=78;
sine[32603]=78;
sine[32604]=78;
sine[32605]=78;
sine[32606]=78;
sine[32607]=78;
sine[32608]=78;
sine[32609]=78;
sine[32610]=78;
sine[32611]=78;
sine[32612]=78;
sine[32613]=78;
sine[32614]=78;
sine[32615]=78;
sine[32616]=78;
sine[32617]=78;
sine[32618]=78;
sine[32619]=78;
sine[32620]=78;
sine[32621]=78;
sine[32622]=78;
sine[32623]=78;
sine[32624]=78;
sine[32625]=78;
sine[32626]=78;
sine[32627]=78;
sine[32628]=78;
sine[32629]=78;
sine[32630]=78;
sine[32631]=78;
sine[32632]=78;
sine[32633]=78;
sine[32634]=78;
sine[32635]=78;
sine[32636]=78;
sine[32637]=78;
sine[32638]=78;
sine[32639]=78;
sine[32640]=78;
sine[32641]=78;
sine[32642]=78;
sine[32643]=78;
sine[32644]=78;
sine[32645]=78;
sine[32646]=78;
sine[32647]=78;
sine[32648]=78;
sine[32649]=78;
sine[32650]=78;
sine[32651]=78;
sine[32652]=78;
sine[32653]=78;
sine[32654]=78;
sine[32655]=78;
sine[32656]=78;
sine[32657]=78;
sine[32658]=78;
sine[32659]=78;
sine[32660]=78;
sine[32661]=78;
sine[32662]=78;
sine[32663]=78;
sine[32664]=78;
sine[32665]=78;
sine[32666]=78;
sine[32667]=78;
sine[32668]=78;
sine[32669]=78;
sine[32670]=78;
sine[32671]=78;
sine[32672]=78;
sine[32673]=78;
sine[32674]=78;
sine[32675]=78;
sine[32676]=78;
sine[32677]=78;
sine[32678]=78;
sine[32679]=78;
sine[32680]=78;
sine[32681]=78;
sine[32682]=78;
sine[32683]=78;
sine[32684]=78;
sine[32685]=78;
sine[32686]=78;
sine[32687]=78;
sine[32688]=78;
sine[32689]=78;
sine[32690]=78;
sine[32691]=78;
sine[32692]=78;
sine[32693]=78;
sine[32694]=78;
sine[32695]=78;
sine[32696]=78;
sine[32697]=78;
sine[32698]=78;
sine[32699]=78;
sine[32700]=78;
sine[32701]=78;
sine[32702]=77;
sine[32703]=77;
sine[32704]=77;
sine[32705]=77;
sine[32706]=77;
sine[32707]=77;
sine[32708]=77;
sine[32709]=77;
sine[32710]=77;
sine[32711]=77;
sine[32712]=77;
sine[32713]=77;
sine[32714]=77;
sine[32715]=77;
sine[32716]=77;
sine[32717]=77;
sine[32718]=77;
sine[32719]=77;
sine[32720]=77;
sine[32721]=77;
sine[32722]=77;
sine[32723]=77;
sine[32724]=77;
sine[32725]=77;
sine[32726]=77;
sine[32727]=77;
sine[32728]=77;
sine[32729]=77;
sine[32730]=77;
sine[32731]=77;
sine[32732]=77;
sine[32733]=77;
sine[32734]=77;
sine[32735]=77;
sine[32736]=77;
sine[32737]=77;
sine[32738]=77;
sine[32739]=77;
sine[32740]=77;
sine[32741]=77;
sine[32742]=77;
sine[32743]=77;
sine[32744]=77;
sine[32745]=77;
sine[32746]=77;
sine[32747]=77;
sine[32748]=77;
sine[32749]=77;
sine[32750]=77;
sine[32751]=77;
sine[32752]=77;
sine[32753]=77;
sine[32754]=77;
sine[32755]=77;
sine[32756]=77;
sine[32757]=77;
sine[32758]=77;
sine[32759]=77;
sine[32760]=77;
sine[32761]=77;
sine[32762]=77;
sine[32763]=77;
sine[32764]=77;
sine[32765]=77;
sine[32766]=77;
sine[32767]=77;
sine[32768]=77;
sine[32769]=77;
sine[32770]=77;
sine[32771]=77;
sine[32772]=77;
sine[32773]=77;
sine[32774]=77;
sine[32775]=77;
sine[32776]=77;
sine[32777]=77;
sine[32778]=77;
sine[32779]=77;
sine[32780]=77;
sine[32781]=77;
sine[32782]=77;
sine[32783]=77;
sine[32784]=77;
sine[32785]=77;
sine[32786]=77;
sine[32787]=77;
sine[32788]=77;
sine[32789]=77;
sine[32790]=77;
sine[32791]=77;
sine[32792]=77;
sine[32793]=77;
sine[32794]=77;
sine[32795]=77;
sine[32796]=77;
sine[32797]=77;
sine[32798]=77;
sine[32799]=77;
sine[32800]=77;
sine[32801]=77;
sine[32802]=77;
sine[32803]=77;
sine[32804]=77;
sine[32805]=77;
sine[32806]=77;
sine[32807]=77;
sine[32808]=77;
sine[32809]=77;
sine[32810]=77;
sine[32811]=77;
sine[32812]=77;
sine[32813]=77;
sine[32814]=77;
sine[32815]=77;
sine[32816]=77;
sine[32817]=77;
sine[32818]=77;
sine[32819]=77;
sine[32820]=77;
sine[32821]=77;
sine[32822]=77;
sine[32823]=77;
sine[32824]=77;
sine[32825]=77;
sine[32826]=76;
sine[32827]=76;
sine[32828]=76;
sine[32829]=76;
sine[32830]=76;
sine[32831]=76;
sine[32832]=76;
sine[32833]=76;
sine[32834]=76;
sine[32835]=76;
sine[32836]=76;
sine[32837]=76;
sine[32838]=76;
sine[32839]=76;
sine[32840]=76;
sine[32841]=76;
sine[32842]=76;
sine[32843]=76;
sine[32844]=76;
sine[32845]=76;
sine[32846]=76;
sine[32847]=76;
sine[32848]=76;
sine[32849]=76;
sine[32850]=76;
sine[32851]=76;
sine[32852]=76;
sine[32853]=76;
sine[32854]=76;
sine[32855]=76;
sine[32856]=76;
sine[32857]=76;
sine[32858]=76;
sine[32859]=76;
sine[32860]=76;
sine[32861]=76;
sine[32862]=76;
sine[32863]=76;
sine[32864]=76;
sine[32865]=76;
sine[32866]=76;
sine[32867]=76;
sine[32868]=76;
sine[32869]=76;
sine[32870]=76;
sine[32871]=76;
sine[32872]=76;
sine[32873]=76;
sine[32874]=76;
sine[32875]=76;
sine[32876]=76;
sine[32877]=76;
sine[32878]=76;
sine[32879]=76;
sine[32880]=76;
sine[32881]=76;
sine[32882]=76;
sine[32883]=76;
sine[32884]=76;
sine[32885]=76;
sine[32886]=76;
sine[32887]=76;
sine[32888]=76;
sine[32889]=76;
sine[32890]=76;
sine[32891]=76;
sine[32892]=76;
sine[32893]=76;
sine[32894]=76;
sine[32895]=76;
sine[32896]=76;
sine[32897]=76;
sine[32898]=76;
sine[32899]=76;
sine[32900]=76;
sine[32901]=76;
sine[32902]=76;
sine[32903]=76;
sine[32904]=76;
sine[32905]=76;
sine[32906]=76;
sine[32907]=76;
sine[32908]=76;
sine[32909]=76;
sine[32910]=76;
sine[32911]=76;
sine[32912]=76;
sine[32913]=76;
sine[32914]=75;
sine[32915]=75;
sine[32916]=75;
sine[32917]=75;
sine[32918]=75;
sine[32919]=75;
sine[32920]=75;
sine[32921]=75;
sine[32922]=75;
sine[32923]=75;
sine[32924]=75;
sine[32925]=75;
sine[32926]=75;
sine[32927]=75;
sine[32928]=75;
sine[32929]=75;
sine[32930]=75;
sine[32931]=75;
sine[32932]=75;
sine[32933]=75;
sine[32934]=75;
sine[32935]=75;
sine[32936]=75;
sine[32937]=75;
sine[32938]=75;
sine[32939]=75;
sine[32940]=75;
sine[32941]=75;
sine[32942]=75;
sine[32943]=75;
sine[32944]=75;
sine[32945]=75;
sine[32946]=75;
sine[32947]=75;
sine[32948]=75;
sine[32949]=75;
sine[32950]=75;
sine[32951]=75;
sine[32952]=75;
sine[32953]=75;
sine[32954]=75;
sine[32955]=75;
sine[32956]=75;
sine[32957]=75;
sine[32958]=75;
sine[32959]=75;
sine[32960]=75;
sine[32961]=75;
sine[32962]=75;
sine[32963]=75;
sine[32964]=75;
sine[32965]=75;
sine[32966]=75;
sine[32967]=75;
sine[32968]=75;
sine[32969]=75;
sine[32970]=75;
sine[32971]=75;
sine[32972]=75;
sine[32973]=75;
sine[32974]=75;
sine[32975]=75;
sine[32976]=75;
sine[32977]=75;
sine[32978]=75;
sine[32979]=75;
sine[32980]=75;
sine[32981]=75;
sine[32982]=75;
sine[32983]=75;
sine[32984]=75;
sine[32985]=75;
sine[32986]=75;
sine[32987]=74;
sine[32988]=74;
sine[32989]=74;
sine[32990]=74;
sine[32991]=74;
sine[32992]=74;
sine[32993]=74;
sine[32994]=74;
sine[32995]=74;
sine[32996]=74;
sine[32997]=74;
sine[32998]=74;
sine[32999]=74;
sine[33000]=74;
sine[33001]=74;
sine[33002]=74;
sine[33003]=74;
sine[33004]=74;
sine[33005]=74;
sine[33006]=74;
sine[33007]=74;
sine[33008]=74;
sine[33009]=74;
sine[33010]=74;
sine[33011]=74;
sine[33012]=74;
sine[33013]=74;
sine[33014]=74;
sine[33015]=74;
sine[33016]=74;
sine[33017]=74;
sine[33018]=74;
sine[33019]=74;
sine[33020]=74;
sine[33021]=74;
sine[33022]=74;
sine[33023]=74;
sine[33024]=74;
sine[33025]=74;
sine[33026]=74;
sine[33027]=74;
sine[33028]=74;
sine[33029]=74;
sine[33030]=74;
sine[33031]=74;
sine[33032]=74;
sine[33033]=74;
sine[33034]=74;
sine[33035]=74;
sine[33036]=74;
sine[33037]=74;
sine[33038]=74;
sine[33039]=74;
sine[33040]=74;
sine[33041]=74;
sine[33042]=74;
sine[33043]=74;
sine[33044]=74;
sine[33045]=74;
sine[33046]=74;
sine[33047]=74;
sine[33048]=74;
sine[33049]=74;
sine[33050]=74;
sine[33051]=73;
sine[33052]=73;
sine[33053]=73;
sine[33054]=73;
sine[33055]=73;
sine[33056]=73;
sine[33057]=73;
sine[33058]=73;
sine[33059]=73;
sine[33060]=73;
sine[33061]=73;
sine[33062]=73;
sine[33063]=73;
sine[33064]=73;
sine[33065]=73;
sine[33066]=73;
sine[33067]=73;
sine[33068]=73;
sine[33069]=73;
sine[33070]=73;
sine[33071]=73;
sine[33072]=73;
sine[33073]=73;
sine[33074]=73;
sine[33075]=73;
sine[33076]=73;
sine[33077]=73;
sine[33078]=73;
sine[33079]=73;
sine[33080]=73;
sine[33081]=73;
sine[33082]=73;
sine[33083]=73;
sine[33084]=73;
sine[33085]=73;
sine[33086]=73;
sine[33087]=73;
sine[33088]=73;
sine[33089]=73;
sine[33090]=73;
sine[33091]=73;
sine[33092]=73;
sine[33093]=73;
sine[33094]=73;
sine[33095]=73;
sine[33096]=73;
sine[33097]=73;
sine[33098]=73;
sine[33099]=73;
sine[33100]=73;
sine[33101]=73;
sine[33102]=73;
sine[33103]=73;
sine[33104]=73;
sine[33105]=73;
sine[33106]=73;
sine[33107]=73;
sine[33108]=72;
sine[33109]=72;
sine[33110]=72;
sine[33111]=72;
sine[33112]=72;
sine[33113]=72;
sine[33114]=72;
sine[33115]=72;
sine[33116]=72;
sine[33117]=72;
sine[33118]=72;
sine[33119]=72;
sine[33120]=72;
sine[33121]=72;
sine[33122]=72;
sine[33123]=72;
sine[33124]=72;
sine[33125]=72;
sine[33126]=72;
sine[33127]=72;
sine[33128]=72;
sine[33129]=72;
sine[33130]=72;
sine[33131]=72;
sine[33132]=72;
sine[33133]=72;
sine[33134]=72;
sine[33135]=72;
sine[33136]=72;
sine[33137]=72;
sine[33138]=72;
sine[33139]=72;
sine[33140]=72;
sine[33141]=72;
sine[33142]=72;
sine[33143]=72;
sine[33144]=72;
sine[33145]=72;
sine[33146]=72;
sine[33147]=72;
sine[33148]=72;
sine[33149]=72;
sine[33150]=72;
sine[33151]=72;
sine[33152]=72;
sine[33153]=72;
sine[33154]=72;
sine[33155]=72;
sine[33156]=72;
sine[33157]=72;
sine[33158]=72;
sine[33159]=72;
sine[33160]=72;
sine[33161]=71;
sine[33162]=71;
sine[33163]=71;
sine[33164]=71;
sine[33165]=71;
sine[33166]=71;
sine[33167]=71;
sine[33168]=71;
sine[33169]=71;
sine[33170]=71;
sine[33171]=71;
sine[33172]=71;
sine[33173]=71;
sine[33174]=71;
sine[33175]=71;
sine[33176]=71;
sine[33177]=71;
sine[33178]=71;
sine[33179]=71;
sine[33180]=71;
sine[33181]=71;
sine[33182]=71;
sine[33183]=71;
sine[33184]=71;
sine[33185]=71;
sine[33186]=71;
sine[33187]=71;
sine[33188]=71;
sine[33189]=71;
sine[33190]=71;
sine[33191]=71;
sine[33192]=71;
sine[33193]=71;
sine[33194]=71;
sine[33195]=71;
sine[33196]=71;
sine[33197]=71;
sine[33198]=71;
sine[33199]=71;
sine[33200]=71;
sine[33201]=71;
sine[33202]=71;
sine[33203]=71;
sine[33204]=71;
sine[33205]=71;
sine[33206]=71;
sine[33207]=71;
sine[33208]=71;
sine[33209]=71;
sine[33210]=70;
sine[33211]=70;
sine[33212]=70;
sine[33213]=70;
sine[33214]=70;
sine[33215]=70;
sine[33216]=70;
sine[33217]=70;
sine[33218]=70;
sine[33219]=70;
sine[33220]=70;
sine[33221]=70;
sine[33222]=70;
sine[33223]=70;
sine[33224]=70;
sine[33225]=70;
sine[33226]=70;
sine[33227]=70;
sine[33228]=70;
sine[33229]=70;
sine[33230]=70;
sine[33231]=70;
sine[33232]=70;
sine[33233]=70;
sine[33234]=70;
sine[33235]=70;
sine[33236]=70;
sine[33237]=70;
sine[33238]=70;
sine[33239]=70;
sine[33240]=70;
sine[33241]=70;
sine[33242]=70;
sine[33243]=70;
sine[33244]=70;
sine[33245]=70;
sine[33246]=70;
sine[33247]=70;
sine[33248]=70;
sine[33249]=70;
sine[33250]=70;
sine[33251]=70;
sine[33252]=70;
sine[33253]=70;
sine[33254]=70;
sine[33255]=69;
sine[33256]=69;
sine[33257]=69;
sine[33258]=69;
sine[33259]=69;
sine[33260]=69;
sine[33261]=69;
sine[33262]=69;
sine[33263]=69;
sine[33264]=69;
sine[33265]=69;
sine[33266]=69;
sine[33267]=69;
sine[33268]=69;
sine[33269]=69;
sine[33270]=69;
sine[33271]=69;
sine[33272]=69;
sine[33273]=69;
sine[33274]=69;
sine[33275]=69;
sine[33276]=69;
sine[33277]=69;
sine[33278]=69;
sine[33279]=69;
sine[33280]=69;
sine[33281]=69;
sine[33282]=69;
sine[33283]=69;
sine[33284]=69;
sine[33285]=69;
sine[33286]=69;
sine[33287]=69;
sine[33288]=69;
sine[33289]=69;
sine[33290]=69;
sine[33291]=69;
sine[33292]=69;
sine[33293]=69;
sine[33294]=69;
sine[33295]=69;
sine[33296]=69;
sine[33297]=69;
sine[33298]=69;
sine[33299]=68;
sine[33300]=68;
sine[33301]=68;
sine[33302]=68;
sine[33303]=68;
sine[33304]=68;
sine[33305]=68;
sine[33306]=68;
sine[33307]=68;
sine[33308]=68;
sine[33309]=68;
sine[33310]=68;
sine[33311]=68;
sine[33312]=68;
sine[33313]=68;
sine[33314]=68;
sine[33315]=68;
sine[33316]=68;
sine[33317]=68;
sine[33318]=68;
sine[33319]=68;
sine[33320]=68;
sine[33321]=68;
sine[33322]=68;
sine[33323]=68;
sine[33324]=68;
sine[33325]=68;
sine[33326]=68;
sine[33327]=68;
sine[33328]=68;
sine[33329]=68;
sine[33330]=68;
sine[33331]=68;
sine[33332]=68;
sine[33333]=68;
sine[33334]=68;
sine[33335]=68;
sine[33336]=68;
sine[33337]=68;
sine[33338]=68;
sine[33339]=68;
sine[33340]=67;
sine[33341]=67;
sine[33342]=67;
sine[33343]=67;
sine[33344]=67;
sine[33345]=67;
sine[33346]=67;
sine[33347]=67;
sine[33348]=67;
sine[33349]=67;
sine[33350]=67;
sine[33351]=67;
sine[33352]=67;
sine[33353]=67;
sine[33354]=67;
sine[33355]=67;
sine[33356]=67;
sine[33357]=67;
sine[33358]=67;
sine[33359]=67;
sine[33360]=67;
sine[33361]=67;
sine[33362]=67;
sine[33363]=67;
sine[33364]=67;
sine[33365]=67;
sine[33366]=67;
sine[33367]=67;
sine[33368]=67;
sine[33369]=67;
sine[33370]=67;
sine[33371]=67;
sine[33372]=67;
sine[33373]=67;
sine[33374]=67;
sine[33375]=67;
sine[33376]=67;
sine[33377]=67;
sine[33378]=67;
sine[33379]=67;
sine[33380]=66;
sine[33381]=66;
sine[33382]=66;
sine[33383]=66;
sine[33384]=66;
sine[33385]=66;
sine[33386]=66;
sine[33387]=66;
sine[33388]=66;
sine[33389]=66;
sine[33390]=66;
sine[33391]=66;
sine[33392]=66;
sine[33393]=66;
sine[33394]=66;
sine[33395]=66;
sine[33396]=66;
sine[33397]=66;
sine[33398]=66;
sine[33399]=66;
sine[33400]=66;
sine[33401]=66;
sine[33402]=66;
sine[33403]=66;
sine[33404]=66;
sine[33405]=66;
sine[33406]=66;
sine[33407]=66;
sine[33408]=66;
sine[33409]=66;
sine[33410]=66;
sine[33411]=66;
sine[33412]=66;
sine[33413]=66;
sine[33414]=66;
sine[33415]=66;
sine[33416]=66;
sine[33417]=66;
sine[33418]=65;
sine[33419]=65;
sine[33420]=65;
sine[33421]=65;
sine[33422]=65;
sine[33423]=65;
sine[33424]=65;
sine[33425]=65;
sine[33426]=65;
sine[33427]=65;
sine[33428]=65;
sine[33429]=65;
sine[33430]=65;
sine[33431]=65;
sine[33432]=65;
sine[33433]=65;
sine[33434]=65;
sine[33435]=65;
sine[33436]=65;
sine[33437]=65;
sine[33438]=65;
sine[33439]=65;
sine[33440]=65;
sine[33441]=65;
sine[33442]=65;
sine[33443]=65;
sine[33444]=65;
sine[33445]=65;
sine[33446]=65;
sine[33447]=65;
sine[33448]=65;
sine[33449]=65;
sine[33450]=65;
sine[33451]=65;
sine[33452]=65;
sine[33453]=65;
sine[33454]=65;
sine[33455]=64;
sine[33456]=64;
sine[33457]=64;
sine[33458]=64;
sine[33459]=64;
sine[33460]=64;
sine[33461]=64;
sine[33462]=64;
sine[33463]=64;
sine[33464]=64;
sine[33465]=64;
sine[33466]=64;
sine[33467]=64;
sine[33468]=64;
sine[33469]=64;
sine[33470]=64;
sine[33471]=64;
sine[33472]=64;
sine[33473]=64;
sine[33474]=64;
sine[33475]=64;
sine[33476]=64;
sine[33477]=64;
sine[33478]=64;
sine[33479]=64;
sine[33480]=64;
sine[33481]=64;
sine[33482]=64;
sine[33483]=64;
sine[33484]=64;
sine[33485]=64;
sine[33486]=64;
sine[33487]=64;
sine[33488]=64;
sine[33489]=64;
sine[33490]=63;
sine[33491]=63;
sine[33492]=63;
sine[33493]=63;
sine[33494]=63;
sine[33495]=63;
sine[33496]=63;
sine[33497]=63;
sine[33498]=63;
sine[33499]=63;
sine[33500]=63;
sine[33501]=63;
sine[33502]=63;
sine[33503]=63;
sine[33504]=63;
sine[33505]=63;
sine[33506]=63;
sine[33507]=63;
sine[33508]=63;
sine[33509]=63;
sine[33510]=63;
sine[33511]=63;
sine[33512]=63;
sine[33513]=63;
sine[33514]=63;
sine[33515]=63;
sine[33516]=63;
sine[33517]=63;
sine[33518]=63;
sine[33519]=63;
sine[33520]=63;
sine[33521]=63;
sine[33522]=63;
sine[33523]=63;
sine[33524]=63;
sine[33525]=62;
sine[33526]=62;
sine[33527]=62;
sine[33528]=62;
sine[33529]=62;
sine[33530]=62;
sine[33531]=62;
sine[33532]=62;
sine[33533]=62;
sine[33534]=62;
sine[33535]=62;
sine[33536]=62;
sine[33537]=62;
sine[33538]=62;
sine[33539]=62;
sine[33540]=62;
sine[33541]=62;
sine[33542]=62;
sine[33543]=62;
sine[33544]=62;
sine[33545]=62;
sine[33546]=62;
sine[33547]=62;
sine[33548]=62;
sine[33549]=62;
sine[33550]=62;
sine[33551]=62;
sine[33552]=62;
sine[33553]=62;
sine[33554]=62;
sine[33555]=62;
sine[33556]=62;
sine[33557]=62;
sine[33558]=61;
sine[33559]=61;
sine[33560]=61;
sine[33561]=61;
sine[33562]=61;
sine[33563]=61;
sine[33564]=61;
sine[33565]=61;
sine[33566]=61;
sine[33567]=61;
sine[33568]=61;
sine[33569]=61;
sine[33570]=61;
sine[33571]=61;
sine[33572]=61;
sine[33573]=61;
sine[33574]=61;
sine[33575]=61;
sine[33576]=61;
sine[33577]=61;
sine[33578]=61;
sine[33579]=61;
sine[33580]=61;
sine[33581]=61;
sine[33582]=61;
sine[33583]=61;
sine[33584]=61;
sine[33585]=61;
sine[33586]=61;
sine[33587]=61;
sine[33588]=61;
sine[33589]=61;
sine[33590]=61;
sine[33591]=60;
sine[33592]=60;
sine[33593]=60;
sine[33594]=60;
sine[33595]=60;
sine[33596]=60;
sine[33597]=60;
sine[33598]=60;
sine[33599]=60;
sine[33600]=60;
sine[33601]=60;
sine[33602]=60;
sine[33603]=60;
sine[33604]=60;
sine[33605]=60;
sine[33606]=60;
sine[33607]=60;
sine[33608]=60;
sine[33609]=60;
sine[33610]=60;
sine[33611]=60;
sine[33612]=60;
sine[33613]=60;
sine[33614]=60;
sine[33615]=60;
sine[33616]=60;
sine[33617]=60;
sine[33618]=60;
sine[33619]=60;
sine[33620]=60;
sine[33621]=60;
sine[33622]=60;
sine[33623]=59;
sine[33624]=59;
sine[33625]=59;
sine[33626]=59;
sine[33627]=59;
sine[33628]=59;
sine[33629]=59;
sine[33630]=59;
sine[33631]=59;
sine[33632]=59;
sine[33633]=59;
sine[33634]=59;
sine[33635]=59;
sine[33636]=59;
sine[33637]=59;
sine[33638]=59;
sine[33639]=59;
sine[33640]=59;
sine[33641]=59;
sine[33642]=59;
sine[33643]=59;
sine[33644]=59;
sine[33645]=59;
sine[33646]=59;
sine[33647]=59;
sine[33648]=59;
sine[33649]=59;
sine[33650]=59;
sine[33651]=59;
sine[33652]=59;
sine[33653]=59;
sine[33654]=58;
sine[33655]=58;
sine[33656]=58;
sine[33657]=58;
sine[33658]=58;
sine[33659]=58;
sine[33660]=58;
sine[33661]=58;
sine[33662]=58;
sine[33663]=58;
sine[33664]=58;
sine[33665]=58;
sine[33666]=58;
sine[33667]=58;
sine[33668]=58;
sine[33669]=58;
sine[33670]=58;
sine[33671]=58;
sine[33672]=58;
sine[33673]=58;
sine[33674]=58;
sine[33675]=58;
sine[33676]=58;
sine[33677]=58;
sine[33678]=58;
sine[33679]=58;
sine[33680]=58;
sine[33681]=58;
sine[33682]=58;
sine[33683]=58;
sine[33684]=57;
sine[33685]=57;
sine[33686]=57;
sine[33687]=57;
sine[33688]=57;
sine[33689]=57;
sine[33690]=57;
sine[33691]=57;
sine[33692]=57;
sine[33693]=57;
sine[33694]=57;
sine[33695]=57;
sine[33696]=57;
sine[33697]=57;
sine[33698]=57;
sine[33699]=57;
sine[33700]=57;
sine[33701]=57;
sine[33702]=57;
sine[33703]=57;
sine[33704]=57;
sine[33705]=57;
sine[33706]=57;
sine[33707]=57;
sine[33708]=57;
sine[33709]=57;
sine[33710]=57;
sine[33711]=57;
sine[33712]=57;
sine[33713]=57;
sine[33714]=56;
sine[33715]=56;
sine[33716]=56;
sine[33717]=56;
sine[33718]=56;
sine[33719]=56;
sine[33720]=56;
sine[33721]=56;
sine[33722]=56;
sine[33723]=56;
sine[33724]=56;
sine[33725]=56;
sine[33726]=56;
sine[33727]=56;
sine[33728]=56;
sine[33729]=56;
sine[33730]=56;
sine[33731]=56;
sine[33732]=56;
sine[33733]=56;
sine[33734]=56;
sine[33735]=56;
sine[33736]=56;
sine[33737]=56;
sine[33738]=56;
sine[33739]=56;
sine[33740]=56;
sine[33741]=56;
sine[33742]=56;
sine[33743]=55;
sine[33744]=55;
sine[33745]=55;
sine[33746]=55;
sine[33747]=55;
sine[33748]=55;
sine[33749]=55;
sine[33750]=55;
sine[33751]=55;
sine[33752]=55;
sine[33753]=55;
sine[33754]=55;
sine[33755]=55;
sine[33756]=55;
sine[33757]=55;
sine[33758]=55;
sine[33759]=55;
sine[33760]=55;
sine[33761]=55;
sine[33762]=55;
sine[33763]=55;
sine[33764]=55;
sine[33765]=55;
sine[33766]=55;
sine[33767]=55;
sine[33768]=55;
sine[33769]=55;
sine[33770]=55;
sine[33771]=55;
sine[33772]=54;
sine[33773]=54;
sine[33774]=54;
sine[33775]=54;
sine[33776]=54;
sine[33777]=54;
sine[33778]=54;
sine[33779]=54;
sine[33780]=54;
sine[33781]=54;
sine[33782]=54;
sine[33783]=54;
sine[33784]=54;
sine[33785]=54;
sine[33786]=54;
sine[33787]=54;
sine[33788]=54;
sine[33789]=54;
sine[33790]=54;
sine[33791]=54;
sine[33792]=54;
sine[33793]=54;
sine[33794]=54;
sine[33795]=54;
sine[33796]=54;
sine[33797]=54;
sine[33798]=54;
sine[33799]=54;
sine[33800]=53;
sine[33801]=53;
sine[33802]=53;
sine[33803]=53;
sine[33804]=53;
sine[33805]=53;
sine[33806]=53;
sine[33807]=53;
sine[33808]=53;
sine[33809]=53;
sine[33810]=53;
sine[33811]=53;
sine[33812]=53;
sine[33813]=53;
sine[33814]=53;
sine[33815]=53;
sine[33816]=53;
sine[33817]=53;
sine[33818]=53;
sine[33819]=53;
sine[33820]=53;
sine[33821]=53;
sine[33822]=53;
sine[33823]=53;
sine[33824]=53;
sine[33825]=53;
sine[33826]=53;
sine[33827]=53;
sine[33828]=52;
sine[33829]=52;
sine[33830]=52;
sine[33831]=52;
sine[33832]=52;
sine[33833]=52;
sine[33834]=52;
sine[33835]=52;
sine[33836]=52;
sine[33837]=52;
sine[33838]=52;
sine[33839]=52;
sine[33840]=52;
sine[33841]=52;
sine[33842]=52;
sine[33843]=52;
sine[33844]=52;
sine[33845]=52;
sine[33846]=52;
sine[33847]=52;
sine[33848]=52;
sine[33849]=52;
sine[33850]=52;
sine[33851]=52;
sine[33852]=52;
sine[33853]=52;
sine[33854]=52;
sine[33855]=51;
sine[33856]=51;
sine[33857]=51;
sine[33858]=51;
sine[33859]=51;
sine[33860]=51;
sine[33861]=51;
sine[33862]=51;
sine[33863]=51;
sine[33864]=51;
sine[33865]=51;
sine[33866]=51;
sine[33867]=51;
sine[33868]=51;
sine[33869]=51;
sine[33870]=51;
sine[33871]=51;
sine[33872]=51;
sine[33873]=51;
sine[33874]=51;
sine[33875]=51;
sine[33876]=51;
sine[33877]=51;
sine[33878]=51;
sine[33879]=51;
sine[33880]=51;
sine[33881]=51;
sine[33882]=50;
sine[33883]=50;
sine[33884]=50;
sine[33885]=50;
sine[33886]=50;
sine[33887]=50;
sine[33888]=50;
sine[33889]=50;
sine[33890]=50;
sine[33891]=50;
sine[33892]=50;
sine[33893]=50;
sine[33894]=50;
sine[33895]=50;
sine[33896]=50;
sine[33897]=50;
sine[33898]=50;
sine[33899]=50;
sine[33900]=50;
sine[33901]=50;
sine[33902]=50;
sine[33903]=50;
sine[33904]=50;
sine[33905]=50;
sine[33906]=50;
sine[33907]=50;
sine[33908]=49;
sine[33909]=49;
sine[33910]=49;
sine[33911]=49;
sine[33912]=49;
sine[33913]=49;
sine[33914]=49;
sine[33915]=49;
sine[33916]=49;
sine[33917]=49;
sine[33918]=49;
sine[33919]=49;
sine[33920]=49;
sine[33921]=49;
sine[33922]=49;
sine[33923]=49;
sine[33924]=49;
sine[33925]=49;
sine[33926]=49;
sine[33927]=49;
sine[33928]=49;
sine[33929]=49;
sine[33930]=49;
sine[33931]=49;
sine[33932]=49;
sine[33933]=49;
sine[33934]=49;
sine[33935]=48;
sine[33936]=48;
sine[33937]=48;
sine[33938]=48;
sine[33939]=48;
sine[33940]=48;
sine[33941]=48;
sine[33942]=48;
sine[33943]=48;
sine[33944]=48;
sine[33945]=48;
sine[33946]=48;
sine[33947]=48;
sine[33948]=48;
sine[33949]=48;
sine[33950]=48;
sine[33951]=48;
sine[33952]=48;
sine[33953]=48;
sine[33954]=48;
sine[33955]=48;
sine[33956]=48;
sine[33957]=48;
sine[33958]=48;
sine[33959]=48;
sine[33960]=47;
sine[33961]=47;
sine[33962]=47;
sine[33963]=47;
sine[33964]=47;
sine[33965]=47;
sine[33966]=47;
sine[33967]=47;
sine[33968]=47;
sine[33969]=47;
sine[33970]=47;
sine[33971]=47;
sine[33972]=47;
sine[33973]=47;
sine[33974]=47;
sine[33975]=47;
sine[33976]=47;
sine[33977]=47;
sine[33978]=47;
sine[33979]=47;
sine[33980]=47;
sine[33981]=47;
sine[33982]=47;
sine[33983]=47;
sine[33984]=47;
sine[33985]=47;
sine[33986]=46;
sine[33987]=46;
sine[33988]=46;
sine[33989]=46;
sine[33990]=46;
sine[33991]=46;
sine[33992]=46;
sine[33993]=46;
sine[33994]=46;
sine[33995]=46;
sine[33996]=46;
sine[33997]=46;
sine[33998]=46;
sine[33999]=46;
sine[34000]=46;
sine[34001]=46;
sine[34002]=46;
sine[34003]=46;
sine[34004]=46;
sine[34005]=46;
sine[34006]=46;
sine[34007]=46;
sine[34008]=46;
sine[34009]=46;
sine[34010]=46;
sine[34011]=45;
sine[34012]=45;
sine[34013]=45;
sine[34014]=45;
sine[34015]=45;
sine[34016]=45;
sine[34017]=45;
sine[34018]=45;
sine[34019]=45;
sine[34020]=45;
sine[34021]=45;
sine[34022]=45;
sine[34023]=45;
sine[34024]=45;
sine[34025]=45;
sine[34026]=45;
sine[34027]=45;
sine[34028]=45;
sine[34029]=45;
sine[34030]=45;
sine[34031]=45;
sine[34032]=45;
sine[34033]=45;
sine[34034]=45;
sine[34035]=45;
sine[34036]=44;
sine[34037]=44;
sine[34038]=44;
sine[34039]=44;
sine[34040]=44;
sine[34041]=44;
sine[34042]=44;
sine[34043]=44;
sine[34044]=44;
sine[34045]=44;
sine[34046]=44;
sine[34047]=44;
sine[34048]=44;
sine[34049]=44;
sine[34050]=44;
sine[34051]=44;
sine[34052]=44;
sine[34053]=44;
sine[34054]=44;
sine[34055]=44;
sine[34056]=44;
sine[34057]=44;
sine[34058]=44;
sine[34059]=44;
sine[34060]=44;
sine[34061]=43;
sine[34062]=43;
sine[34063]=43;
sine[34064]=43;
sine[34065]=43;
sine[34066]=43;
sine[34067]=43;
sine[34068]=43;
sine[34069]=43;
sine[34070]=43;
sine[34071]=43;
sine[34072]=43;
sine[34073]=43;
sine[34074]=43;
sine[34075]=43;
sine[34076]=43;
sine[34077]=43;
sine[34078]=43;
sine[34079]=43;
sine[34080]=43;
sine[34081]=43;
sine[34082]=43;
sine[34083]=43;
sine[34084]=43;
sine[34085]=42;
sine[34086]=42;
sine[34087]=42;
sine[34088]=42;
sine[34089]=42;
sine[34090]=42;
sine[34091]=42;
sine[34092]=42;
sine[34093]=42;
sine[34094]=42;
sine[34095]=42;
sine[34096]=42;
sine[34097]=42;
sine[34098]=42;
sine[34099]=42;
sine[34100]=42;
sine[34101]=42;
sine[34102]=42;
sine[34103]=42;
sine[34104]=42;
sine[34105]=42;
sine[34106]=42;
sine[34107]=42;
sine[34108]=42;
sine[34109]=41;
sine[34110]=41;
sine[34111]=41;
sine[34112]=41;
sine[34113]=41;
sine[34114]=41;
sine[34115]=41;
sine[34116]=41;
sine[34117]=41;
sine[34118]=41;
sine[34119]=41;
sine[34120]=41;
sine[34121]=41;
sine[34122]=41;
sine[34123]=41;
sine[34124]=41;
sine[34125]=41;
sine[34126]=41;
sine[34127]=41;
sine[34128]=41;
sine[34129]=41;
sine[34130]=41;
sine[34131]=41;
sine[34132]=41;
sine[34133]=40;
sine[34134]=40;
sine[34135]=40;
sine[34136]=40;
sine[34137]=40;
sine[34138]=40;
sine[34139]=40;
sine[34140]=40;
sine[34141]=40;
sine[34142]=40;
sine[34143]=40;
sine[34144]=40;
sine[34145]=40;
sine[34146]=40;
sine[34147]=40;
sine[34148]=40;
sine[34149]=40;
sine[34150]=40;
sine[34151]=40;
sine[34152]=40;
sine[34153]=40;
sine[34154]=40;
sine[34155]=40;
sine[34156]=40;
sine[34157]=39;
sine[34158]=39;
sine[34159]=39;
sine[34160]=39;
sine[34161]=39;
sine[34162]=39;
sine[34163]=39;
sine[34164]=39;
sine[34165]=39;
sine[34166]=39;
sine[34167]=39;
sine[34168]=39;
sine[34169]=39;
sine[34170]=39;
sine[34171]=39;
sine[34172]=39;
sine[34173]=39;
sine[34174]=39;
sine[34175]=39;
sine[34176]=39;
sine[34177]=39;
sine[34178]=39;
sine[34179]=39;
sine[34180]=38;
sine[34181]=38;
sine[34182]=38;
sine[34183]=38;
sine[34184]=38;
sine[34185]=38;
sine[34186]=38;
sine[34187]=38;
sine[34188]=38;
sine[34189]=38;
sine[34190]=38;
sine[34191]=38;
sine[34192]=38;
sine[34193]=38;
sine[34194]=38;
sine[34195]=38;
sine[34196]=38;
sine[34197]=38;
sine[34198]=38;
sine[34199]=38;
sine[34200]=38;
sine[34201]=38;
sine[34202]=38;
sine[34203]=38;
sine[34204]=37;
sine[34205]=37;
sine[34206]=37;
sine[34207]=37;
sine[34208]=37;
sine[34209]=37;
sine[34210]=37;
sine[34211]=37;
sine[34212]=37;
sine[34213]=37;
sine[34214]=37;
sine[34215]=37;
sine[34216]=37;
sine[34217]=37;
sine[34218]=37;
sine[34219]=37;
sine[34220]=37;
sine[34221]=37;
sine[34222]=37;
sine[34223]=37;
sine[34224]=37;
sine[34225]=37;
sine[34226]=37;
sine[34227]=36;
sine[34228]=36;
sine[34229]=36;
sine[34230]=36;
sine[34231]=36;
sine[34232]=36;
sine[34233]=36;
sine[34234]=36;
sine[34235]=36;
sine[34236]=36;
sine[34237]=36;
sine[34238]=36;
sine[34239]=36;
sine[34240]=36;
sine[34241]=36;
sine[34242]=36;
sine[34243]=36;
sine[34244]=36;
sine[34245]=36;
sine[34246]=36;
sine[34247]=36;
sine[34248]=36;
sine[34249]=36;
sine[34250]=35;
sine[34251]=35;
sine[34252]=35;
sine[34253]=35;
sine[34254]=35;
sine[34255]=35;
sine[34256]=35;
sine[34257]=35;
sine[34258]=35;
sine[34259]=35;
sine[34260]=35;
sine[34261]=35;
sine[34262]=35;
sine[34263]=35;
sine[34264]=35;
sine[34265]=35;
sine[34266]=35;
sine[34267]=35;
sine[34268]=35;
sine[34269]=35;
sine[34270]=35;
sine[34271]=35;
sine[34272]=35;
sine[34273]=34;
sine[34274]=34;
sine[34275]=34;
sine[34276]=34;
sine[34277]=34;
sine[34278]=34;
sine[34279]=34;
sine[34280]=34;
sine[34281]=34;
sine[34282]=34;
sine[34283]=34;
sine[34284]=34;
sine[34285]=34;
sine[34286]=34;
sine[34287]=34;
sine[34288]=34;
sine[34289]=34;
sine[34290]=34;
sine[34291]=34;
sine[34292]=34;
sine[34293]=34;
sine[34294]=34;
sine[34295]=33;
sine[34296]=33;
sine[34297]=33;
sine[34298]=33;
sine[34299]=33;
sine[34300]=33;
sine[34301]=33;
sine[34302]=33;
sine[34303]=33;
sine[34304]=33;
sine[34305]=33;
sine[34306]=33;
sine[34307]=33;
sine[34308]=33;
sine[34309]=33;
sine[34310]=33;
sine[34311]=33;
sine[34312]=33;
sine[34313]=33;
sine[34314]=33;
sine[34315]=33;
sine[34316]=33;
sine[34317]=33;
sine[34318]=32;
sine[34319]=32;
sine[34320]=32;
sine[34321]=32;
sine[34322]=32;
sine[34323]=32;
sine[34324]=32;
sine[34325]=32;
sine[34326]=32;
sine[34327]=32;
sine[34328]=32;
sine[34329]=32;
sine[34330]=32;
sine[34331]=32;
sine[34332]=32;
sine[34333]=32;
sine[34334]=32;
sine[34335]=32;
sine[34336]=32;
sine[34337]=32;
sine[34338]=32;
sine[34339]=32;
sine[34340]=31;
sine[34341]=31;
sine[34342]=31;
sine[34343]=31;
sine[34344]=31;
sine[34345]=31;
sine[34346]=31;
sine[34347]=31;
sine[34348]=31;
sine[34349]=31;
sine[34350]=31;
sine[34351]=31;
sine[34352]=31;
sine[34353]=31;
sine[34354]=31;
sine[34355]=31;
sine[34356]=31;
sine[34357]=31;
sine[34358]=31;
sine[34359]=31;
sine[34360]=31;
sine[34361]=31;
sine[34362]=30;
sine[34363]=30;
sine[34364]=30;
sine[34365]=30;
sine[34366]=30;
sine[34367]=30;
sine[34368]=30;
sine[34369]=30;
sine[34370]=30;
sine[34371]=30;
sine[34372]=30;
sine[34373]=30;
sine[34374]=30;
sine[34375]=30;
sine[34376]=30;
sine[34377]=30;
sine[34378]=30;
sine[34379]=30;
sine[34380]=30;
sine[34381]=30;
sine[34382]=30;
sine[34383]=30;
sine[34384]=29;
sine[34385]=29;
sine[34386]=29;
sine[34387]=29;
sine[34388]=29;
sine[34389]=29;
sine[34390]=29;
sine[34391]=29;
sine[34392]=29;
sine[34393]=29;
sine[34394]=29;
sine[34395]=29;
sine[34396]=29;
sine[34397]=29;
sine[34398]=29;
sine[34399]=29;
sine[34400]=29;
sine[34401]=29;
sine[34402]=29;
sine[34403]=29;
sine[34404]=29;
sine[34405]=29;
sine[34406]=28;
sine[34407]=28;
sine[34408]=28;
sine[34409]=28;
sine[34410]=28;
sine[34411]=28;
sine[34412]=28;
sine[34413]=28;
sine[34414]=28;
sine[34415]=28;
sine[34416]=28;
sine[34417]=28;
sine[34418]=28;
sine[34419]=28;
sine[34420]=28;
sine[34421]=28;
sine[34422]=28;
sine[34423]=28;
sine[34424]=28;
sine[34425]=28;
sine[34426]=28;
sine[34427]=28;
sine[34428]=27;
sine[34429]=27;
sine[34430]=27;
sine[34431]=27;
sine[34432]=27;
sine[34433]=27;
sine[34434]=27;
sine[34435]=27;
sine[34436]=27;
sine[34437]=27;
sine[34438]=27;
sine[34439]=27;
sine[34440]=27;
sine[34441]=27;
sine[34442]=27;
sine[34443]=27;
sine[34444]=27;
sine[34445]=27;
sine[34446]=27;
sine[34447]=27;
sine[34448]=27;
sine[34449]=27;
sine[34450]=26;
sine[34451]=26;
sine[34452]=26;
sine[34453]=26;
sine[34454]=26;
sine[34455]=26;
sine[34456]=26;
sine[34457]=26;
sine[34458]=26;
sine[34459]=26;
sine[34460]=26;
sine[34461]=26;
sine[34462]=26;
sine[34463]=26;
sine[34464]=26;
sine[34465]=26;
sine[34466]=26;
sine[34467]=26;
sine[34468]=26;
sine[34469]=26;
sine[34470]=26;
sine[34471]=25;
sine[34472]=25;
sine[34473]=25;
sine[34474]=25;
sine[34475]=25;
sine[34476]=25;
sine[34477]=25;
sine[34478]=25;
sine[34479]=25;
sine[34480]=25;
sine[34481]=25;
sine[34482]=25;
sine[34483]=25;
sine[34484]=25;
sine[34485]=25;
sine[34486]=25;
sine[34487]=25;
sine[34488]=25;
sine[34489]=25;
sine[34490]=25;
sine[34491]=25;
sine[34492]=25;
sine[34493]=24;
sine[34494]=24;
sine[34495]=24;
sine[34496]=24;
sine[34497]=24;
sine[34498]=24;
sine[34499]=24;
sine[34500]=24;
sine[34501]=24;
sine[34502]=24;
sine[34503]=24;
sine[34504]=24;
sine[34505]=24;
sine[34506]=24;
sine[34507]=24;
sine[34508]=24;
sine[34509]=24;
sine[34510]=24;
sine[34511]=24;
sine[34512]=24;
sine[34513]=24;
sine[34514]=23;
sine[34515]=23;
sine[34516]=23;
sine[34517]=23;
sine[34518]=23;
sine[34519]=23;
sine[34520]=23;
sine[34521]=23;
sine[34522]=23;
sine[34523]=23;
sine[34524]=23;
sine[34525]=23;
sine[34526]=23;
sine[34527]=23;
sine[34528]=23;
sine[34529]=23;
sine[34530]=23;
sine[34531]=23;
sine[34532]=23;
sine[34533]=23;
sine[34534]=23;
sine[34535]=23;
sine[34536]=22;
sine[34537]=22;
sine[34538]=22;
sine[34539]=22;
sine[34540]=22;
sine[34541]=22;
sine[34542]=22;
sine[34543]=22;
sine[34544]=22;
sine[34545]=22;
sine[34546]=22;
sine[34547]=22;
sine[34548]=22;
sine[34549]=22;
sine[34550]=22;
sine[34551]=22;
sine[34552]=22;
sine[34553]=22;
sine[34554]=22;
sine[34555]=22;
sine[34556]=22;
sine[34557]=21;
sine[34558]=21;
sine[34559]=21;
sine[34560]=21;
sine[34561]=21;
sine[34562]=21;
sine[34563]=21;
sine[34564]=21;
sine[34565]=21;
sine[34566]=21;
sine[34567]=21;
sine[34568]=21;
sine[34569]=21;
sine[34570]=21;
sine[34571]=21;
sine[34572]=21;
sine[34573]=21;
sine[34574]=21;
sine[34575]=21;
sine[34576]=21;
sine[34577]=21;
sine[34578]=20;
sine[34579]=20;
sine[34580]=20;
sine[34581]=20;
sine[34582]=20;
sine[34583]=20;
sine[34584]=20;
sine[34585]=20;
sine[34586]=20;
sine[34587]=20;
sine[34588]=20;
sine[34589]=20;
sine[34590]=20;
sine[34591]=20;
sine[34592]=20;
sine[34593]=20;
sine[34594]=20;
sine[34595]=20;
sine[34596]=20;
sine[34597]=20;
sine[34598]=20;
sine[34599]=19;
sine[34600]=19;
sine[34601]=19;
sine[34602]=19;
sine[34603]=19;
sine[34604]=19;
sine[34605]=19;
sine[34606]=19;
sine[34607]=19;
sine[34608]=19;
sine[34609]=19;
sine[34610]=19;
sine[34611]=19;
sine[34612]=19;
sine[34613]=19;
sine[34614]=19;
sine[34615]=19;
sine[34616]=19;
sine[34617]=19;
sine[34618]=19;
sine[34619]=19;
sine[34620]=18;
sine[34621]=18;
sine[34622]=18;
sine[34623]=18;
sine[34624]=18;
sine[34625]=18;
sine[34626]=18;
sine[34627]=18;
sine[34628]=18;
sine[34629]=18;
sine[34630]=18;
sine[34631]=18;
sine[34632]=18;
sine[34633]=18;
sine[34634]=18;
sine[34635]=18;
sine[34636]=18;
sine[34637]=18;
sine[34638]=18;
sine[34639]=18;
sine[34640]=18;
sine[34641]=17;
sine[34642]=17;
sine[34643]=17;
sine[34644]=17;
sine[34645]=17;
sine[34646]=17;
sine[34647]=17;
sine[34648]=17;
sine[34649]=17;
sine[34650]=17;
sine[34651]=17;
sine[34652]=17;
sine[34653]=17;
sine[34654]=17;
sine[34655]=17;
sine[34656]=17;
sine[34657]=17;
sine[34658]=17;
sine[34659]=17;
sine[34660]=17;
sine[34661]=17;
sine[34662]=16;
sine[34663]=16;
sine[34664]=16;
sine[34665]=16;
sine[34666]=16;
sine[34667]=16;
sine[34668]=16;
sine[34669]=16;
sine[34670]=16;
sine[34671]=16;
sine[34672]=16;
sine[34673]=16;
sine[34674]=16;
sine[34675]=16;
sine[34676]=16;
sine[34677]=16;
sine[34678]=16;
sine[34679]=16;
sine[34680]=16;
sine[34681]=16;
sine[34682]=16;
sine[34683]=15;
sine[34684]=15;
sine[34685]=15;
sine[34686]=15;
sine[34687]=15;
sine[34688]=15;
sine[34689]=15;
sine[34690]=15;
sine[34691]=15;
sine[34692]=15;
sine[34693]=15;
sine[34694]=15;
sine[34695]=15;
sine[34696]=15;
sine[34697]=15;
sine[34698]=15;
sine[34699]=15;
sine[34700]=15;
sine[34701]=15;
sine[34702]=15;
sine[34703]=14;
sine[34704]=14;
sine[34705]=14;
sine[34706]=14;
sine[34707]=14;
sine[34708]=14;
sine[34709]=14;
sine[34710]=14;
sine[34711]=14;
sine[34712]=14;
sine[34713]=14;
sine[34714]=14;
sine[34715]=14;
sine[34716]=14;
sine[34717]=14;
sine[34718]=14;
sine[34719]=14;
sine[34720]=14;
sine[34721]=14;
sine[34722]=14;
sine[34723]=14;
sine[34724]=13;
sine[34725]=13;
sine[34726]=13;
sine[34727]=13;
sine[34728]=13;
sine[34729]=13;
sine[34730]=13;
sine[34731]=13;
sine[34732]=13;
sine[34733]=13;
sine[34734]=13;
sine[34735]=13;
sine[34736]=13;
sine[34737]=13;
sine[34738]=13;
sine[34739]=13;
sine[34740]=13;
sine[34741]=13;
sine[34742]=13;
sine[34743]=13;
sine[34744]=13;
sine[34745]=12;
sine[34746]=12;
sine[34747]=12;
sine[34748]=12;
sine[34749]=12;
sine[34750]=12;
sine[34751]=12;
sine[34752]=12;
sine[34753]=12;
sine[34754]=12;
sine[34755]=12;
sine[34756]=12;
sine[34757]=12;
sine[34758]=12;
sine[34759]=12;
sine[34760]=12;
sine[34761]=12;
sine[34762]=12;
sine[34763]=12;
sine[34764]=12;
sine[34765]=11;
sine[34766]=11;
sine[34767]=11;
sine[34768]=11;
sine[34769]=11;
sine[34770]=11;
sine[34771]=11;
sine[34772]=11;
sine[34773]=11;
sine[34774]=11;
sine[34775]=11;
sine[34776]=11;
sine[34777]=11;
sine[34778]=11;
sine[34779]=11;
sine[34780]=11;
sine[34781]=11;
sine[34782]=11;
sine[34783]=11;
sine[34784]=11;
sine[34785]=11;
sine[34786]=10;
sine[34787]=10;
sine[34788]=10;
sine[34789]=10;
sine[34790]=10;
sine[34791]=10;
sine[34792]=10;
sine[34793]=10;
sine[34794]=10;
sine[34795]=10;
sine[34796]=10;
sine[34797]=10;
sine[34798]=10;
sine[34799]=10;
sine[34800]=10;
sine[34801]=10;
sine[34802]=10;
sine[34803]=10;
sine[34804]=10;
sine[34805]=10;
sine[34806]=9;
sine[34807]=9;
sine[34808]=9;
sine[34809]=9;
sine[34810]=9;
sine[34811]=9;
sine[34812]=9;
sine[34813]=9;
sine[34814]=9;
sine[34815]=9;
sine[34816]=9;
sine[34817]=9;
sine[34818]=9;
sine[34819]=9;
sine[34820]=9;
sine[34821]=9;
sine[34822]=9;
sine[34823]=9;
sine[34824]=9;
sine[34825]=9;
sine[34826]=9;
sine[34827]=8;
sine[34828]=8;
sine[34829]=8;
sine[34830]=8;
sine[34831]=8;
sine[34832]=8;
sine[34833]=8;
sine[34834]=8;
sine[34835]=8;
sine[34836]=8;
sine[34837]=8;
sine[34838]=8;
sine[34839]=8;
sine[34840]=8;
sine[34841]=8;
sine[34842]=8;
sine[34843]=8;
sine[34844]=8;
sine[34845]=8;
sine[34846]=8;
sine[34847]=7;
sine[34848]=7;
sine[34849]=7;
sine[34850]=7;
sine[34851]=7;
sine[34852]=7;
sine[34853]=7;
sine[34854]=7;
sine[34855]=7;
sine[34856]=7;
sine[34857]=7;
sine[34858]=7;
sine[34859]=7;
sine[34860]=7;
sine[34861]=7;
sine[34862]=7;
sine[34863]=7;
sine[34864]=7;
sine[34865]=7;
sine[34866]=7;
sine[34867]=7;
sine[34868]=6;
sine[34869]=6;
sine[34870]=6;
sine[34871]=6;
sine[34872]=6;
sine[34873]=6;
sine[34874]=6;
sine[34875]=6;
sine[34876]=6;
sine[34877]=6;
sine[34878]=6;
sine[34879]=6;
sine[34880]=6;
sine[34881]=6;
sine[34882]=6;
sine[34883]=6;
sine[34884]=6;
sine[34885]=6;
sine[34886]=6;
sine[34887]=6;
sine[34888]=5;
sine[34889]=5;
sine[34890]=5;
sine[34891]=5;
sine[34892]=5;
sine[34893]=5;
sine[34894]=5;
sine[34895]=5;
sine[34896]=5;
sine[34897]=5;
sine[34898]=5;
sine[34899]=5;
sine[34900]=5;
sine[34901]=5;
sine[34902]=5;
sine[34903]=5;
sine[34904]=5;
sine[34905]=5;
sine[34906]=5;
sine[34907]=5;
sine[34908]=5;
sine[34909]=4;
sine[34910]=4;
sine[34911]=4;
sine[34912]=4;
sine[34913]=4;
sine[34914]=4;
sine[34915]=4;
sine[34916]=4;
sine[34917]=4;
sine[34918]=4;
sine[34919]=4;
sine[34920]=4;
sine[34921]=4;
sine[34922]=4;
sine[34923]=4;
sine[34924]=4;
sine[34925]=4;
sine[34926]=4;
sine[34927]=4;
sine[34928]=4;
sine[34929]=3;
sine[34930]=3;
sine[34931]=3;
sine[34932]=3;
sine[34933]=3;
sine[34934]=3;
sine[34935]=3;
sine[34936]=3;
sine[34937]=3;
sine[34938]=3;
sine[34939]=3;
sine[34940]=3;
sine[34941]=3;
sine[34942]=3;
sine[34943]=3;
sine[34944]=3;
sine[34945]=3;
sine[34946]=3;
sine[34947]=3;
sine[34948]=3;
sine[34949]=3;
sine[34950]=2;
sine[34951]=2;
sine[34952]=2;
sine[34953]=2;
sine[34954]=2;
sine[34955]=2;
sine[34956]=2;
sine[34957]=2;
sine[34958]=2;
sine[34959]=2;
sine[34960]=2;
sine[34961]=2;
sine[34962]=2;
sine[34963]=2;
sine[34964]=2;
sine[34965]=2;
sine[34966]=2;
sine[34967]=2;
sine[34968]=2;
sine[34969]=2;
sine[34970]=1;
sine[34971]=1;
sine[34972]=1;
sine[34973]=1;
sine[34974]=1;
sine[34975]=1;
sine[34976]=1;
sine[34977]=1;
sine[34978]=1;
sine[34979]=1;
sine[34980]=1;
sine[34981]=1;
sine[34982]=1;
sine[34983]=1;
sine[34984]=1;
sine[34985]=1;
sine[34986]=1;
sine[34987]=1;
sine[34988]=1;
sine[34989]=1;
sine[34990]=0;
sine[34991]=0;
sine[34992]=0;
sine[34993]=0;
sine[34994]=0;
sine[34995]=0;
sine[34996]=0;
sine[34997]=0;
sine[34998]=0;
sine[34999]=0;
sine[35000]=0;
sine[35001]=0;
sine[35002]=0;
sine[35003]=0;
sine[35004]=0;
sine[35005]=0;
sine[35006]=0;
sine[35007]=0;
sine[35008]=0;
sine[35009]=0;
sine[35010]=0;
sine[35011]=-1;
sine[35012]=-1;
sine[35013]=-1;
sine[35014]=-1;
sine[35015]=-1;
sine[35016]=-1;
sine[35017]=-1;
sine[35018]=-1;
sine[35019]=-1;
sine[35020]=-1;
sine[35021]=-1;
sine[35022]=-1;
sine[35023]=-1;
sine[35024]=-1;
sine[35025]=-1;
sine[35026]=-1;
sine[35027]=-1;
sine[35028]=-1;
sine[35029]=-1;
sine[35030]=-1;
sine[35031]=-2;
sine[35032]=-2;
sine[35033]=-2;
sine[35034]=-2;
sine[35035]=-2;
sine[35036]=-2;
sine[35037]=-2;
sine[35038]=-2;
sine[35039]=-2;
sine[35040]=-2;
sine[35041]=-2;
sine[35042]=-2;
sine[35043]=-2;
sine[35044]=-2;
sine[35045]=-2;
sine[35046]=-2;
sine[35047]=-2;
sine[35048]=-2;
sine[35049]=-2;
sine[35050]=-2;
sine[35051]=-3;
sine[35052]=-3;
sine[35053]=-3;
sine[35054]=-3;
sine[35055]=-3;
sine[35056]=-3;
sine[35057]=-3;
sine[35058]=-3;
sine[35059]=-3;
sine[35060]=-3;
sine[35061]=-3;
sine[35062]=-3;
sine[35063]=-3;
sine[35064]=-3;
sine[35065]=-3;
sine[35066]=-3;
sine[35067]=-3;
sine[35068]=-3;
sine[35069]=-3;
sine[35070]=-3;
sine[35071]=-3;
sine[35072]=-4;
sine[35073]=-4;
sine[35074]=-4;
sine[35075]=-4;
sine[35076]=-4;
sine[35077]=-4;
sine[35078]=-4;
sine[35079]=-4;
sine[35080]=-4;
sine[35081]=-4;
sine[35082]=-4;
sine[35083]=-4;
sine[35084]=-4;
sine[35085]=-4;
sine[35086]=-4;
sine[35087]=-4;
sine[35088]=-4;
sine[35089]=-4;
sine[35090]=-4;
sine[35091]=-4;
sine[35092]=-5;
sine[35093]=-5;
sine[35094]=-5;
sine[35095]=-5;
sine[35096]=-5;
sine[35097]=-5;
sine[35098]=-5;
sine[35099]=-5;
sine[35100]=-5;
sine[35101]=-5;
sine[35102]=-5;
sine[35103]=-5;
sine[35104]=-5;
sine[35105]=-5;
sine[35106]=-5;
sine[35107]=-5;
sine[35108]=-5;
sine[35109]=-5;
sine[35110]=-5;
sine[35111]=-5;
sine[35112]=-5;
sine[35113]=-6;
sine[35114]=-6;
sine[35115]=-6;
sine[35116]=-6;
sine[35117]=-6;
sine[35118]=-6;
sine[35119]=-6;
sine[35120]=-6;
sine[35121]=-6;
sine[35122]=-6;
sine[35123]=-6;
sine[35124]=-6;
sine[35125]=-6;
sine[35126]=-6;
sine[35127]=-6;
sine[35128]=-6;
sine[35129]=-6;
sine[35130]=-6;
sine[35131]=-6;
sine[35132]=-6;
sine[35133]=-7;
sine[35134]=-7;
sine[35135]=-7;
sine[35136]=-7;
sine[35137]=-7;
sine[35138]=-7;
sine[35139]=-7;
sine[35140]=-7;
sine[35141]=-7;
sine[35142]=-7;
sine[35143]=-7;
sine[35144]=-7;
sine[35145]=-7;
sine[35146]=-7;
sine[35147]=-7;
sine[35148]=-7;
sine[35149]=-7;
sine[35150]=-7;
sine[35151]=-7;
sine[35152]=-7;
sine[35153]=-7;
sine[35154]=-8;
sine[35155]=-8;
sine[35156]=-8;
sine[35157]=-8;
sine[35158]=-8;
sine[35159]=-8;
sine[35160]=-8;
sine[35161]=-8;
sine[35162]=-8;
sine[35163]=-8;
sine[35164]=-8;
sine[35165]=-8;
sine[35166]=-8;
sine[35167]=-8;
sine[35168]=-8;
sine[35169]=-8;
sine[35170]=-8;
sine[35171]=-8;
sine[35172]=-8;
sine[35173]=-8;
sine[35174]=-9;
sine[35175]=-9;
sine[35176]=-9;
sine[35177]=-9;
sine[35178]=-9;
sine[35179]=-9;
sine[35180]=-9;
sine[35181]=-9;
sine[35182]=-9;
sine[35183]=-9;
sine[35184]=-9;
sine[35185]=-9;
sine[35186]=-9;
sine[35187]=-9;
sine[35188]=-9;
sine[35189]=-9;
sine[35190]=-9;
sine[35191]=-9;
sine[35192]=-9;
sine[35193]=-9;
sine[35194]=-9;
sine[35195]=-10;
sine[35196]=-10;
sine[35197]=-10;
sine[35198]=-10;
sine[35199]=-10;
sine[35200]=-10;
sine[35201]=-10;
sine[35202]=-10;
sine[35203]=-10;
sine[35204]=-10;
sine[35205]=-10;
sine[35206]=-10;
sine[35207]=-10;
sine[35208]=-10;
sine[35209]=-10;
sine[35210]=-10;
sine[35211]=-10;
sine[35212]=-10;
sine[35213]=-10;
sine[35214]=-10;
sine[35215]=-11;
sine[35216]=-11;
sine[35217]=-11;
sine[35218]=-11;
sine[35219]=-11;
sine[35220]=-11;
sine[35221]=-11;
sine[35222]=-11;
sine[35223]=-11;
sine[35224]=-11;
sine[35225]=-11;
sine[35226]=-11;
sine[35227]=-11;
sine[35228]=-11;
sine[35229]=-11;
sine[35230]=-11;
sine[35231]=-11;
sine[35232]=-11;
sine[35233]=-11;
sine[35234]=-11;
sine[35235]=-11;
sine[35236]=-12;
sine[35237]=-12;
sine[35238]=-12;
sine[35239]=-12;
sine[35240]=-12;
sine[35241]=-12;
sine[35242]=-12;
sine[35243]=-12;
sine[35244]=-12;
sine[35245]=-12;
sine[35246]=-12;
sine[35247]=-12;
sine[35248]=-12;
sine[35249]=-12;
sine[35250]=-12;
sine[35251]=-12;
sine[35252]=-12;
sine[35253]=-12;
sine[35254]=-12;
sine[35255]=-12;
sine[35256]=-13;
sine[35257]=-13;
sine[35258]=-13;
sine[35259]=-13;
sine[35260]=-13;
sine[35261]=-13;
sine[35262]=-13;
sine[35263]=-13;
sine[35264]=-13;
sine[35265]=-13;
sine[35266]=-13;
sine[35267]=-13;
sine[35268]=-13;
sine[35269]=-13;
sine[35270]=-13;
sine[35271]=-13;
sine[35272]=-13;
sine[35273]=-13;
sine[35274]=-13;
sine[35275]=-13;
sine[35276]=-13;
sine[35277]=-14;
sine[35278]=-14;
sine[35279]=-14;
sine[35280]=-14;
sine[35281]=-14;
sine[35282]=-14;
sine[35283]=-14;
sine[35284]=-14;
sine[35285]=-14;
sine[35286]=-14;
sine[35287]=-14;
sine[35288]=-14;
sine[35289]=-14;
sine[35290]=-14;
sine[35291]=-14;
sine[35292]=-14;
sine[35293]=-14;
sine[35294]=-14;
sine[35295]=-14;
sine[35296]=-14;
sine[35297]=-14;
sine[35298]=-15;
sine[35299]=-15;
sine[35300]=-15;
sine[35301]=-15;
sine[35302]=-15;
sine[35303]=-15;
sine[35304]=-15;
sine[35305]=-15;
sine[35306]=-15;
sine[35307]=-15;
sine[35308]=-15;
sine[35309]=-15;
sine[35310]=-15;
sine[35311]=-15;
sine[35312]=-15;
sine[35313]=-15;
sine[35314]=-15;
sine[35315]=-15;
sine[35316]=-15;
sine[35317]=-15;
sine[35318]=-16;
sine[35319]=-16;
sine[35320]=-16;
sine[35321]=-16;
sine[35322]=-16;
sine[35323]=-16;
sine[35324]=-16;
sine[35325]=-16;
sine[35326]=-16;
sine[35327]=-16;
sine[35328]=-16;
sine[35329]=-16;
sine[35330]=-16;
sine[35331]=-16;
sine[35332]=-16;
sine[35333]=-16;
sine[35334]=-16;
sine[35335]=-16;
sine[35336]=-16;
sine[35337]=-16;
sine[35338]=-16;
sine[35339]=-17;
sine[35340]=-17;
sine[35341]=-17;
sine[35342]=-17;
sine[35343]=-17;
sine[35344]=-17;
sine[35345]=-17;
sine[35346]=-17;
sine[35347]=-17;
sine[35348]=-17;
sine[35349]=-17;
sine[35350]=-17;
sine[35351]=-17;
sine[35352]=-17;
sine[35353]=-17;
sine[35354]=-17;
sine[35355]=-17;
sine[35356]=-17;
sine[35357]=-17;
sine[35358]=-17;
sine[35359]=-17;
sine[35360]=-18;
sine[35361]=-18;
sine[35362]=-18;
sine[35363]=-18;
sine[35364]=-18;
sine[35365]=-18;
sine[35366]=-18;
sine[35367]=-18;
sine[35368]=-18;
sine[35369]=-18;
sine[35370]=-18;
sine[35371]=-18;
sine[35372]=-18;
sine[35373]=-18;
sine[35374]=-18;
sine[35375]=-18;
sine[35376]=-18;
sine[35377]=-18;
sine[35378]=-18;
sine[35379]=-18;
sine[35380]=-18;
sine[35381]=-19;
sine[35382]=-19;
sine[35383]=-19;
sine[35384]=-19;
sine[35385]=-19;
sine[35386]=-19;
sine[35387]=-19;
sine[35388]=-19;
sine[35389]=-19;
sine[35390]=-19;
sine[35391]=-19;
sine[35392]=-19;
sine[35393]=-19;
sine[35394]=-19;
sine[35395]=-19;
sine[35396]=-19;
sine[35397]=-19;
sine[35398]=-19;
sine[35399]=-19;
sine[35400]=-19;
sine[35401]=-19;
sine[35402]=-20;
sine[35403]=-20;
sine[35404]=-20;
sine[35405]=-20;
sine[35406]=-20;
sine[35407]=-20;
sine[35408]=-20;
sine[35409]=-20;
sine[35410]=-20;
sine[35411]=-20;
sine[35412]=-20;
sine[35413]=-20;
sine[35414]=-20;
sine[35415]=-20;
sine[35416]=-20;
sine[35417]=-20;
sine[35418]=-20;
sine[35419]=-20;
sine[35420]=-20;
sine[35421]=-20;
sine[35422]=-20;
sine[35423]=-21;
sine[35424]=-21;
sine[35425]=-21;
sine[35426]=-21;
sine[35427]=-21;
sine[35428]=-21;
sine[35429]=-21;
sine[35430]=-21;
sine[35431]=-21;
sine[35432]=-21;
sine[35433]=-21;
sine[35434]=-21;
sine[35435]=-21;
sine[35436]=-21;
sine[35437]=-21;
sine[35438]=-21;
sine[35439]=-21;
sine[35440]=-21;
sine[35441]=-21;
sine[35442]=-21;
sine[35443]=-21;
sine[35444]=-22;
sine[35445]=-22;
sine[35446]=-22;
sine[35447]=-22;
sine[35448]=-22;
sine[35449]=-22;
sine[35450]=-22;
sine[35451]=-22;
sine[35452]=-22;
sine[35453]=-22;
sine[35454]=-22;
sine[35455]=-22;
sine[35456]=-22;
sine[35457]=-22;
sine[35458]=-22;
sine[35459]=-22;
sine[35460]=-22;
sine[35461]=-22;
sine[35462]=-22;
sine[35463]=-22;
sine[35464]=-22;
sine[35465]=-23;
sine[35466]=-23;
sine[35467]=-23;
sine[35468]=-23;
sine[35469]=-23;
sine[35470]=-23;
sine[35471]=-23;
sine[35472]=-23;
sine[35473]=-23;
sine[35474]=-23;
sine[35475]=-23;
sine[35476]=-23;
sine[35477]=-23;
sine[35478]=-23;
sine[35479]=-23;
sine[35480]=-23;
sine[35481]=-23;
sine[35482]=-23;
sine[35483]=-23;
sine[35484]=-23;
sine[35485]=-23;
sine[35486]=-23;
sine[35487]=-24;
sine[35488]=-24;
sine[35489]=-24;
sine[35490]=-24;
sine[35491]=-24;
sine[35492]=-24;
sine[35493]=-24;
sine[35494]=-24;
sine[35495]=-24;
sine[35496]=-24;
sine[35497]=-24;
sine[35498]=-24;
sine[35499]=-24;
sine[35500]=-24;
sine[35501]=-24;
sine[35502]=-24;
sine[35503]=-24;
sine[35504]=-24;
sine[35505]=-24;
sine[35506]=-24;
sine[35507]=-24;
sine[35508]=-25;
sine[35509]=-25;
sine[35510]=-25;
sine[35511]=-25;
sine[35512]=-25;
sine[35513]=-25;
sine[35514]=-25;
sine[35515]=-25;
sine[35516]=-25;
sine[35517]=-25;
sine[35518]=-25;
sine[35519]=-25;
sine[35520]=-25;
sine[35521]=-25;
sine[35522]=-25;
sine[35523]=-25;
sine[35524]=-25;
sine[35525]=-25;
sine[35526]=-25;
sine[35527]=-25;
sine[35528]=-25;
sine[35529]=-25;
sine[35530]=-26;
sine[35531]=-26;
sine[35532]=-26;
sine[35533]=-26;
sine[35534]=-26;
sine[35535]=-26;
sine[35536]=-26;
sine[35537]=-26;
sine[35538]=-26;
sine[35539]=-26;
sine[35540]=-26;
sine[35541]=-26;
sine[35542]=-26;
sine[35543]=-26;
sine[35544]=-26;
sine[35545]=-26;
sine[35546]=-26;
sine[35547]=-26;
sine[35548]=-26;
sine[35549]=-26;
sine[35550]=-26;
sine[35551]=-27;
sine[35552]=-27;
sine[35553]=-27;
sine[35554]=-27;
sine[35555]=-27;
sine[35556]=-27;
sine[35557]=-27;
sine[35558]=-27;
sine[35559]=-27;
sine[35560]=-27;
sine[35561]=-27;
sine[35562]=-27;
sine[35563]=-27;
sine[35564]=-27;
sine[35565]=-27;
sine[35566]=-27;
sine[35567]=-27;
sine[35568]=-27;
sine[35569]=-27;
sine[35570]=-27;
sine[35571]=-27;
sine[35572]=-27;
sine[35573]=-28;
sine[35574]=-28;
sine[35575]=-28;
sine[35576]=-28;
sine[35577]=-28;
sine[35578]=-28;
sine[35579]=-28;
sine[35580]=-28;
sine[35581]=-28;
sine[35582]=-28;
sine[35583]=-28;
sine[35584]=-28;
sine[35585]=-28;
sine[35586]=-28;
sine[35587]=-28;
sine[35588]=-28;
sine[35589]=-28;
sine[35590]=-28;
sine[35591]=-28;
sine[35592]=-28;
sine[35593]=-28;
sine[35594]=-28;
sine[35595]=-29;
sine[35596]=-29;
sine[35597]=-29;
sine[35598]=-29;
sine[35599]=-29;
sine[35600]=-29;
sine[35601]=-29;
sine[35602]=-29;
sine[35603]=-29;
sine[35604]=-29;
sine[35605]=-29;
sine[35606]=-29;
sine[35607]=-29;
sine[35608]=-29;
sine[35609]=-29;
sine[35610]=-29;
sine[35611]=-29;
sine[35612]=-29;
sine[35613]=-29;
sine[35614]=-29;
sine[35615]=-29;
sine[35616]=-29;
sine[35617]=-30;
sine[35618]=-30;
sine[35619]=-30;
sine[35620]=-30;
sine[35621]=-30;
sine[35622]=-30;
sine[35623]=-30;
sine[35624]=-30;
sine[35625]=-30;
sine[35626]=-30;
sine[35627]=-30;
sine[35628]=-30;
sine[35629]=-30;
sine[35630]=-30;
sine[35631]=-30;
sine[35632]=-30;
sine[35633]=-30;
sine[35634]=-30;
sine[35635]=-30;
sine[35636]=-30;
sine[35637]=-30;
sine[35638]=-30;
sine[35639]=-31;
sine[35640]=-31;
sine[35641]=-31;
sine[35642]=-31;
sine[35643]=-31;
sine[35644]=-31;
sine[35645]=-31;
sine[35646]=-31;
sine[35647]=-31;
sine[35648]=-31;
sine[35649]=-31;
sine[35650]=-31;
sine[35651]=-31;
sine[35652]=-31;
sine[35653]=-31;
sine[35654]=-31;
sine[35655]=-31;
sine[35656]=-31;
sine[35657]=-31;
sine[35658]=-31;
sine[35659]=-31;
sine[35660]=-31;
sine[35661]=-32;
sine[35662]=-32;
sine[35663]=-32;
sine[35664]=-32;
sine[35665]=-32;
sine[35666]=-32;
sine[35667]=-32;
sine[35668]=-32;
sine[35669]=-32;
sine[35670]=-32;
sine[35671]=-32;
sine[35672]=-32;
sine[35673]=-32;
sine[35674]=-32;
sine[35675]=-32;
sine[35676]=-32;
sine[35677]=-32;
sine[35678]=-32;
sine[35679]=-32;
sine[35680]=-32;
sine[35681]=-32;
sine[35682]=-32;
sine[35683]=-33;
sine[35684]=-33;
sine[35685]=-33;
sine[35686]=-33;
sine[35687]=-33;
sine[35688]=-33;
sine[35689]=-33;
sine[35690]=-33;
sine[35691]=-33;
sine[35692]=-33;
sine[35693]=-33;
sine[35694]=-33;
sine[35695]=-33;
sine[35696]=-33;
sine[35697]=-33;
sine[35698]=-33;
sine[35699]=-33;
sine[35700]=-33;
sine[35701]=-33;
sine[35702]=-33;
sine[35703]=-33;
sine[35704]=-33;
sine[35705]=-33;
sine[35706]=-34;
sine[35707]=-34;
sine[35708]=-34;
sine[35709]=-34;
sine[35710]=-34;
sine[35711]=-34;
sine[35712]=-34;
sine[35713]=-34;
sine[35714]=-34;
sine[35715]=-34;
sine[35716]=-34;
sine[35717]=-34;
sine[35718]=-34;
sine[35719]=-34;
sine[35720]=-34;
sine[35721]=-34;
sine[35722]=-34;
sine[35723]=-34;
sine[35724]=-34;
sine[35725]=-34;
sine[35726]=-34;
sine[35727]=-34;
sine[35728]=-35;
sine[35729]=-35;
sine[35730]=-35;
sine[35731]=-35;
sine[35732]=-35;
sine[35733]=-35;
sine[35734]=-35;
sine[35735]=-35;
sine[35736]=-35;
sine[35737]=-35;
sine[35738]=-35;
sine[35739]=-35;
sine[35740]=-35;
sine[35741]=-35;
sine[35742]=-35;
sine[35743]=-35;
sine[35744]=-35;
sine[35745]=-35;
sine[35746]=-35;
sine[35747]=-35;
sine[35748]=-35;
sine[35749]=-35;
sine[35750]=-35;
sine[35751]=-36;
sine[35752]=-36;
sine[35753]=-36;
sine[35754]=-36;
sine[35755]=-36;
sine[35756]=-36;
sine[35757]=-36;
sine[35758]=-36;
sine[35759]=-36;
sine[35760]=-36;
sine[35761]=-36;
sine[35762]=-36;
sine[35763]=-36;
sine[35764]=-36;
sine[35765]=-36;
sine[35766]=-36;
sine[35767]=-36;
sine[35768]=-36;
sine[35769]=-36;
sine[35770]=-36;
sine[35771]=-36;
sine[35772]=-36;
sine[35773]=-36;
sine[35774]=-37;
sine[35775]=-37;
sine[35776]=-37;
sine[35777]=-37;
sine[35778]=-37;
sine[35779]=-37;
sine[35780]=-37;
sine[35781]=-37;
sine[35782]=-37;
sine[35783]=-37;
sine[35784]=-37;
sine[35785]=-37;
sine[35786]=-37;
sine[35787]=-37;
sine[35788]=-37;
sine[35789]=-37;
sine[35790]=-37;
sine[35791]=-37;
sine[35792]=-37;
sine[35793]=-37;
sine[35794]=-37;
sine[35795]=-37;
sine[35796]=-37;
sine[35797]=-38;
sine[35798]=-38;
sine[35799]=-38;
sine[35800]=-38;
sine[35801]=-38;
sine[35802]=-38;
sine[35803]=-38;
sine[35804]=-38;
sine[35805]=-38;
sine[35806]=-38;
sine[35807]=-38;
sine[35808]=-38;
sine[35809]=-38;
sine[35810]=-38;
sine[35811]=-38;
sine[35812]=-38;
sine[35813]=-38;
sine[35814]=-38;
sine[35815]=-38;
sine[35816]=-38;
sine[35817]=-38;
sine[35818]=-38;
sine[35819]=-38;
sine[35820]=-38;
sine[35821]=-39;
sine[35822]=-39;
sine[35823]=-39;
sine[35824]=-39;
sine[35825]=-39;
sine[35826]=-39;
sine[35827]=-39;
sine[35828]=-39;
sine[35829]=-39;
sine[35830]=-39;
sine[35831]=-39;
sine[35832]=-39;
sine[35833]=-39;
sine[35834]=-39;
sine[35835]=-39;
sine[35836]=-39;
sine[35837]=-39;
sine[35838]=-39;
sine[35839]=-39;
sine[35840]=-39;
sine[35841]=-39;
sine[35842]=-39;
sine[35843]=-39;
sine[35844]=-40;
sine[35845]=-40;
sine[35846]=-40;
sine[35847]=-40;
sine[35848]=-40;
sine[35849]=-40;
sine[35850]=-40;
sine[35851]=-40;
sine[35852]=-40;
sine[35853]=-40;
sine[35854]=-40;
sine[35855]=-40;
sine[35856]=-40;
sine[35857]=-40;
sine[35858]=-40;
sine[35859]=-40;
sine[35860]=-40;
sine[35861]=-40;
sine[35862]=-40;
sine[35863]=-40;
sine[35864]=-40;
sine[35865]=-40;
sine[35866]=-40;
sine[35867]=-40;
sine[35868]=-41;
sine[35869]=-41;
sine[35870]=-41;
sine[35871]=-41;
sine[35872]=-41;
sine[35873]=-41;
sine[35874]=-41;
sine[35875]=-41;
sine[35876]=-41;
sine[35877]=-41;
sine[35878]=-41;
sine[35879]=-41;
sine[35880]=-41;
sine[35881]=-41;
sine[35882]=-41;
sine[35883]=-41;
sine[35884]=-41;
sine[35885]=-41;
sine[35886]=-41;
sine[35887]=-41;
sine[35888]=-41;
sine[35889]=-41;
sine[35890]=-41;
sine[35891]=-41;
sine[35892]=-42;
sine[35893]=-42;
sine[35894]=-42;
sine[35895]=-42;
sine[35896]=-42;
sine[35897]=-42;
sine[35898]=-42;
sine[35899]=-42;
sine[35900]=-42;
sine[35901]=-42;
sine[35902]=-42;
sine[35903]=-42;
sine[35904]=-42;
sine[35905]=-42;
sine[35906]=-42;
sine[35907]=-42;
sine[35908]=-42;
sine[35909]=-42;
sine[35910]=-42;
sine[35911]=-42;
sine[35912]=-42;
sine[35913]=-42;
sine[35914]=-42;
sine[35915]=-42;
sine[35916]=-43;
sine[35917]=-43;
sine[35918]=-43;
sine[35919]=-43;
sine[35920]=-43;
sine[35921]=-43;
sine[35922]=-43;
sine[35923]=-43;
sine[35924]=-43;
sine[35925]=-43;
sine[35926]=-43;
sine[35927]=-43;
sine[35928]=-43;
sine[35929]=-43;
sine[35930]=-43;
sine[35931]=-43;
sine[35932]=-43;
sine[35933]=-43;
sine[35934]=-43;
sine[35935]=-43;
sine[35936]=-43;
sine[35937]=-43;
sine[35938]=-43;
sine[35939]=-43;
sine[35940]=-44;
sine[35941]=-44;
sine[35942]=-44;
sine[35943]=-44;
sine[35944]=-44;
sine[35945]=-44;
sine[35946]=-44;
sine[35947]=-44;
sine[35948]=-44;
sine[35949]=-44;
sine[35950]=-44;
sine[35951]=-44;
sine[35952]=-44;
sine[35953]=-44;
sine[35954]=-44;
sine[35955]=-44;
sine[35956]=-44;
sine[35957]=-44;
sine[35958]=-44;
sine[35959]=-44;
sine[35960]=-44;
sine[35961]=-44;
sine[35962]=-44;
sine[35963]=-44;
sine[35964]=-44;
sine[35965]=-45;
sine[35966]=-45;
sine[35967]=-45;
sine[35968]=-45;
sine[35969]=-45;
sine[35970]=-45;
sine[35971]=-45;
sine[35972]=-45;
sine[35973]=-45;
sine[35974]=-45;
sine[35975]=-45;
sine[35976]=-45;
sine[35977]=-45;
sine[35978]=-45;
sine[35979]=-45;
sine[35980]=-45;
sine[35981]=-45;
sine[35982]=-45;
sine[35983]=-45;
sine[35984]=-45;
sine[35985]=-45;
sine[35986]=-45;
sine[35987]=-45;
sine[35988]=-45;
sine[35989]=-45;
sine[35990]=-46;
sine[35991]=-46;
sine[35992]=-46;
sine[35993]=-46;
sine[35994]=-46;
sine[35995]=-46;
sine[35996]=-46;
sine[35997]=-46;
sine[35998]=-46;
sine[35999]=-46;
sine[36000]=-46;
sine[36001]=-46;
sine[36002]=-46;
sine[36003]=-46;
sine[36004]=-46;
sine[36005]=-46;
sine[36006]=-46;
sine[36007]=-46;
sine[36008]=-46;
sine[36009]=-46;
sine[36010]=-46;
sine[36011]=-46;
sine[36012]=-46;
sine[36013]=-46;
sine[36014]=-46;
sine[36015]=-47;
sine[36016]=-47;
sine[36017]=-47;
sine[36018]=-47;
sine[36019]=-47;
sine[36020]=-47;
sine[36021]=-47;
sine[36022]=-47;
sine[36023]=-47;
sine[36024]=-47;
sine[36025]=-47;
sine[36026]=-47;
sine[36027]=-47;
sine[36028]=-47;
sine[36029]=-47;
sine[36030]=-47;
sine[36031]=-47;
sine[36032]=-47;
sine[36033]=-47;
sine[36034]=-47;
sine[36035]=-47;
sine[36036]=-47;
sine[36037]=-47;
sine[36038]=-47;
sine[36039]=-47;
sine[36040]=-47;
sine[36041]=-48;
sine[36042]=-48;
sine[36043]=-48;
sine[36044]=-48;
sine[36045]=-48;
sine[36046]=-48;
sine[36047]=-48;
sine[36048]=-48;
sine[36049]=-48;
sine[36050]=-48;
sine[36051]=-48;
sine[36052]=-48;
sine[36053]=-48;
sine[36054]=-48;
sine[36055]=-48;
sine[36056]=-48;
sine[36057]=-48;
sine[36058]=-48;
sine[36059]=-48;
sine[36060]=-48;
sine[36061]=-48;
sine[36062]=-48;
sine[36063]=-48;
sine[36064]=-48;
sine[36065]=-48;
sine[36066]=-49;
sine[36067]=-49;
sine[36068]=-49;
sine[36069]=-49;
sine[36070]=-49;
sine[36071]=-49;
sine[36072]=-49;
sine[36073]=-49;
sine[36074]=-49;
sine[36075]=-49;
sine[36076]=-49;
sine[36077]=-49;
sine[36078]=-49;
sine[36079]=-49;
sine[36080]=-49;
sine[36081]=-49;
sine[36082]=-49;
sine[36083]=-49;
sine[36084]=-49;
sine[36085]=-49;
sine[36086]=-49;
sine[36087]=-49;
sine[36088]=-49;
sine[36089]=-49;
sine[36090]=-49;
sine[36091]=-49;
sine[36092]=-49;
sine[36093]=-50;
sine[36094]=-50;
sine[36095]=-50;
sine[36096]=-50;
sine[36097]=-50;
sine[36098]=-50;
sine[36099]=-50;
sine[36100]=-50;
sine[36101]=-50;
sine[36102]=-50;
sine[36103]=-50;
sine[36104]=-50;
sine[36105]=-50;
sine[36106]=-50;
sine[36107]=-50;
sine[36108]=-50;
sine[36109]=-50;
sine[36110]=-50;
sine[36111]=-50;
sine[36112]=-50;
sine[36113]=-50;
sine[36114]=-50;
sine[36115]=-50;
sine[36116]=-50;
sine[36117]=-50;
sine[36118]=-50;
sine[36119]=-51;
sine[36120]=-51;
sine[36121]=-51;
sine[36122]=-51;
sine[36123]=-51;
sine[36124]=-51;
sine[36125]=-51;
sine[36126]=-51;
sine[36127]=-51;
sine[36128]=-51;
sine[36129]=-51;
sine[36130]=-51;
sine[36131]=-51;
sine[36132]=-51;
sine[36133]=-51;
sine[36134]=-51;
sine[36135]=-51;
sine[36136]=-51;
sine[36137]=-51;
sine[36138]=-51;
sine[36139]=-51;
sine[36140]=-51;
sine[36141]=-51;
sine[36142]=-51;
sine[36143]=-51;
sine[36144]=-51;
sine[36145]=-51;
sine[36146]=-52;
sine[36147]=-52;
sine[36148]=-52;
sine[36149]=-52;
sine[36150]=-52;
sine[36151]=-52;
sine[36152]=-52;
sine[36153]=-52;
sine[36154]=-52;
sine[36155]=-52;
sine[36156]=-52;
sine[36157]=-52;
sine[36158]=-52;
sine[36159]=-52;
sine[36160]=-52;
sine[36161]=-52;
sine[36162]=-52;
sine[36163]=-52;
sine[36164]=-52;
sine[36165]=-52;
sine[36166]=-52;
sine[36167]=-52;
sine[36168]=-52;
sine[36169]=-52;
sine[36170]=-52;
sine[36171]=-52;
sine[36172]=-52;
sine[36173]=-53;
sine[36174]=-53;
sine[36175]=-53;
sine[36176]=-53;
sine[36177]=-53;
sine[36178]=-53;
sine[36179]=-53;
sine[36180]=-53;
sine[36181]=-53;
sine[36182]=-53;
sine[36183]=-53;
sine[36184]=-53;
sine[36185]=-53;
sine[36186]=-53;
sine[36187]=-53;
sine[36188]=-53;
sine[36189]=-53;
sine[36190]=-53;
sine[36191]=-53;
sine[36192]=-53;
sine[36193]=-53;
sine[36194]=-53;
sine[36195]=-53;
sine[36196]=-53;
sine[36197]=-53;
sine[36198]=-53;
sine[36199]=-53;
sine[36200]=-53;
sine[36201]=-54;
sine[36202]=-54;
sine[36203]=-54;
sine[36204]=-54;
sine[36205]=-54;
sine[36206]=-54;
sine[36207]=-54;
sine[36208]=-54;
sine[36209]=-54;
sine[36210]=-54;
sine[36211]=-54;
sine[36212]=-54;
sine[36213]=-54;
sine[36214]=-54;
sine[36215]=-54;
sine[36216]=-54;
sine[36217]=-54;
sine[36218]=-54;
sine[36219]=-54;
sine[36220]=-54;
sine[36221]=-54;
sine[36222]=-54;
sine[36223]=-54;
sine[36224]=-54;
sine[36225]=-54;
sine[36226]=-54;
sine[36227]=-54;
sine[36228]=-54;
sine[36229]=-55;
sine[36230]=-55;
sine[36231]=-55;
sine[36232]=-55;
sine[36233]=-55;
sine[36234]=-55;
sine[36235]=-55;
sine[36236]=-55;
sine[36237]=-55;
sine[36238]=-55;
sine[36239]=-55;
sine[36240]=-55;
sine[36241]=-55;
sine[36242]=-55;
sine[36243]=-55;
sine[36244]=-55;
sine[36245]=-55;
sine[36246]=-55;
sine[36247]=-55;
sine[36248]=-55;
sine[36249]=-55;
sine[36250]=-55;
sine[36251]=-55;
sine[36252]=-55;
sine[36253]=-55;
sine[36254]=-55;
sine[36255]=-55;
sine[36256]=-55;
sine[36257]=-55;
sine[36258]=-56;
sine[36259]=-56;
sine[36260]=-56;
sine[36261]=-56;
sine[36262]=-56;
sine[36263]=-56;
sine[36264]=-56;
sine[36265]=-56;
sine[36266]=-56;
sine[36267]=-56;
sine[36268]=-56;
sine[36269]=-56;
sine[36270]=-56;
sine[36271]=-56;
sine[36272]=-56;
sine[36273]=-56;
sine[36274]=-56;
sine[36275]=-56;
sine[36276]=-56;
sine[36277]=-56;
sine[36278]=-56;
sine[36279]=-56;
sine[36280]=-56;
sine[36281]=-56;
sine[36282]=-56;
sine[36283]=-56;
sine[36284]=-56;
sine[36285]=-56;
sine[36286]=-56;
sine[36287]=-57;
sine[36288]=-57;
sine[36289]=-57;
sine[36290]=-57;
sine[36291]=-57;
sine[36292]=-57;
sine[36293]=-57;
sine[36294]=-57;
sine[36295]=-57;
sine[36296]=-57;
sine[36297]=-57;
sine[36298]=-57;
sine[36299]=-57;
sine[36300]=-57;
sine[36301]=-57;
sine[36302]=-57;
sine[36303]=-57;
sine[36304]=-57;
sine[36305]=-57;
sine[36306]=-57;
sine[36307]=-57;
sine[36308]=-57;
sine[36309]=-57;
sine[36310]=-57;
sine[36311]=-57;
sine[36312]=-57;
sine[36313]=-57;
sine[36314]=-57;
sine[36315]=-57;
sine[36316]=-57;
sine[36317]=-58;
sine[36318]=-58;
sine[36319]=-58;
sine[36320]=-58;
sine[36321]=-58;
sine[36322]=-58;
sine[36323]=-58;
sine[36324]=-58;
sine[36325]=-58;
sine[36326]=-58;
sine[36327]=-58;
sine[36328]=-58;
sine[36329]=-58;
sine[36330]=-58;
sine[36331]=-58;
sine[36332]=-58;
sine[36333]=-58;
sine[36334]=-58;
sine[36335]=-58;
sine[36336]=-58;
sine[36337]=-58;
sine[36338]=-58;
sine[36339]=-58;
sine[36340]=-58;
sine[36341]=-58;
sine[36342]=-58;
sine[36343]=-58;
sine[36344]=-58;
sine[36345]=-58;
sine[36346]=-58;
sine[36347]=-59;
sine[36348]=-59;
sine[36349]=-59;
sine[36350]=-59;
sine[36351]=-59;
sine[36352]=-59;
sine[36353]=-59;
sine[36354]=-59;
sine[36355]=-59;
sine[36356]=-59;
sine[36357]=-59;
sine[36358]=-59;
sine[36359]=-59;
sine[36360]=-59;
sine[36361]=-59;
sine[36362]=-59;
sine[36363]=-59;
sine[36364]=-59;
sine[36365]=-59;
sine[36366]=-59;
sine[36367]=-59;
sine[36368]=-59;
sine[36369]=-59;
sine[36370]=-59;
sine[36371]=-59;
sine[36372]=-59;
sine[36373]=-59;
sine[36374]=-59;
sine[36375]=-59;
sine[36376]=-59;
sine[36377]=-59;
sine[36378]=-60;
sine[36379]=-60;
sine[36380]=-60;
sine[36381]=-60;
sine[36382]=-60;
sine[36383]=-60;
sine[36384]=-60;
sine[36385]=-60;
sine[36386]=-60;
sine[36387]=-60;
sine[36388]=-60;
sine[36389]=-60;
sine[36390]=-60;
sine[36391]=-60;
sine[36392]=-60;
sine[36393]=-60;
sine[36394]=-60;
sine[36395]=-60;
sine[36396]=-60;
sine[36397]=-60;
sine[36398]=-60;
sine[36399]=-60;
sine[36400]=-60;
sine[36401]=-60;
sine[36402]=-60;
sine[36403]=-60;
sine[36404]=-60;
sine[36405]=-60;
sine[36406]=-60;
sine[36407]=-60;
sine[36408]=-60;
sine[36409]=-60;
sine[36410]=-61;
sine[36411]=-61;
sine[36412]=-61;
sine[36413]=-61;
sine[36414]=-61;
sine[36415]=-61;
sine[36416]=-61;
sine[36417]=-61;
sine[36418]=-61;
sine[36419]=-61;
sine[36420]=-61;
sine[36421]=-61;
sine[36422]=-61;
sine[36423]=-61;
sine[36424]=-61;
sine[36425]=-61;
sine[36426]=-61;
sine[36427]=-61;
sine[36428]=-61;
sine[36429]=-61;
sine[36430]=-61;
sine[36431]=-61;
sine[36432]=-61;
sine[36433]=-61;
sine[36434]=-61;
sine[36435]=-61;
sine[36436]=-61;
sine[36437]=-61;
sine[36438]=-61;
sine[36439]=-61;
sine[36440]=-61;
sine[36441]=-61;
sine[36442]=-61;
sine[36443]=-62;
sine[36444]=-62;
sine[36445]=-62;
sine[36446]=-62;
sine[36447]=-62;
sine[36448]=-62;
sine[36449]=-62;
sine[36450]=-62;
sine[36451]=-62;
sine[36452]=-62;
sine[36453]=-62;
sine[36454]=-62;
sine[36455]=-62;
sine[36456]=-62;
sine[36457]=-62;
sine[36458]=-62;
sine[36459]=-62;
sine[36460]=-62;
sine[36461]=-62;
sine[36462]=-62;
sine[36463]=-62;
sine[36464]=-62;
sine[36465]=-62;
sine[36466]=-62;
sine[36467]=-62;
sine[36468]=-62;
sine[36469]=-62;
sine[36470]=-62;
sine[36471]=-62;
sine[36472]=-62;
sine[36473]=-62;
sine[36474]=-62;
sine[36475]=-62;
sine[36476]=-63;
sine[36477]=-63;
sine[36478]=-63;
sine[36479]=-63;
sine[36480]=-63;
sine[36481]=-63;
sine[36482]=-63;
sine[36483]=-63;
sine[36484]=-63;
sine[36485]=-63;
sine[36486]=-63;
sine[36487]=-63;
sine[36488]=-63;
sine[36489]=-63;
sine[36490]=-63;
sine[36491]=-63;
sine[36492]=-63;
sine[36493]=-63;
sine[36494]=-63;
sine[36495]=-63;
sine[36496]=-63;
sine[36497]=-63;
sine[36498]=-63;
sine[36499]=-63;
sine[36500]=-63;
sine[36501]=-63;
sine[36502]=-63;
sine[36503]=-63;
sine[36504]=-63;
sine[36505]=-63;
sine[36506]=-63;
sine[36507]=-63;
sine[36508]=-63;
sine[36509]=-63;
sine[36510]=-63;
sine[36511]=-64;
sine[36512]=-64;
sine[36513]=-64;
sine[36514]=-64;
sine[36515]=-64;
sine[36516]=-64;
sine[36517]=-64;
sine[36518]=-64;
sine[36519]=-64;
sine[36520]=-64;
sine[36521]=-64;
sine[36522]=-64;
sine[36523]=-64;
sine[36524]=-64;
sine[36525]=-64;
sine[36526]=-64;
sine[36527]=-64;
sine[36528]=-64;
sine[36529]=-64;
sine[36530]=-64;
sine[36531]=-64;
sine[36532]=-64;
sine[36533]=-64;
sine[36534]=-64;
sine[36535]=-64;
sine[36536]=-64;
sine[36537]=-64;
sine[36538]=-64;
sine[36539]=-64;
sine[36540]=-64;
sine[36541]=-64;
sine[36542]=-64;
sine[36543]=-64;
sine[36544]=-64;
sine[36545]=-64;
sine[36546]=-65;
sine[36547]=-65;
sine[36548]=-65;
sine[36549]=-65;
sine[36550]=-65;
sine[36551]=-65;
sine[36552]=-65;
sine[36553]=-65;
sine[36554]=-65;
sine[36555]=-65;
sine[36556]=-65;
sine[36557]=-65;
sine[36558]=-65;
sine[36559]=-65;
sine[36560]=-65;
sine[36561]=-65;
sine[36562]=-65;
sine[36563]=-65;
sine[36564]=-65;
sine[36565]=-65;
sine[36566]=-65;
sine[36567]=-65;
sine[36568]=-65;
sine[36569]=-65;
sine[36570]=-65;
sine[36571]=-65;
sine[36572]=-65;
sine[36573]=-65;
sine[36574]=-65;
sine[36575]=-65;
sine[36576]=-65;
sine[36577]=-65;
sine[36578]=-65;
sine[36579]=-65;
sine[36580]=-65;
sine[36581]=-65;
sine[36582]=-65;
sine[36583]=-66;
sine[36584]=-66;
sine[36585]=-66;
sine[36586]=-66;
sine[36587]=-66;
sine[36588]=-66;
sine[36589]=-66;
sine[36590]=-66;
sine[36591]=-66;
sine[36592]=-66;
sine[36593]=-66;
sine[36594]=-66;
sine[36595]=-66;
sine[36596]=-66;
sine[36597]=-66;
sine[36598]=-66;
sine[36599]=-66;
sine[36600]=-66;
sine[36601]=-66;
sine[36602]=-66;
sine[36603]=-66;
sine[36604]=-66;
sine[36605]=-66;
sine[36606]=-66;
sine[36607]=-66;
sine[36608]=-66;
sine[36609]=-66;
sine[36610]=-66;
sine[36611]=-66;
sine[36612]=-66;
sine[36613]=-66;
sine[36614]=-66;
sine[36615]=-66;
sine[36616]=-66;
sine[36617]=-66;
sine[36618]=-66;
sine[36619]=-66;
sine[36620]=-66;
sine[36621]=-67;
sine[36622]=-67;
sine[36623]=-67;
sine[36624]=-67;
sine[36625]=-67;
sine[36626]=-67;
sine[36627]=-67;
sine[36628]=-67;
sine[36629]=-67;
sine[36630]=-67;
sine[36631]=-67;
sine[36632]=-67;
sine[36633]=-67;
sine[36634]=-67;
sine[36635]=-67;
sine[36636]=-67;
sine[36637]=-67;
sine[36638]=-67;
sine[36639]=-67;
sine[36640]=-67;
sine[36641]=-67;
sine[36642]=-67;
sine[36643]=-67;
sine[36644]=-67;
sine[36645]=-67;
sine[36646]=-67;
sine[36647]=-67;
sine[36648]=-67;
sine[36649]=-67;
sine[36650]=-67;
sine[36651]=-67;
sine[36652]=-67;
sine[36653]=-67;
sine[36654]=-67;
sine[36655]=-67;
sine[36656]=-67;
sine[36657]=-67;
sine[36658]=-67;
sine[36659]=-67;
sine[36660]=-67;
sine[36661]=-68;
sine[36662]=-68;
sine[36663]=-68;
sine[36664]=-68;
sine[36665]=-68;
sine[36666]=-68;
sine[36667]=-68;
sine[36668]=-68;
sine[36669]=-68;
sine[36670]=-68;
sine[36671]=-68;
sine[36672]=-68;
sine[36673]=-68;
sine[36674]=-68;
sine[36675]=-68;
sine[36676]=-68;
sine[36677]=-68;
sine[36678]=-68;
sine[36679]=-68;
sine[36680]=-68;
sine[36681]=-68;
sine[36682]=-68;
sine[36683]=-68;
sine[36684]=-68;
sine[36685]=-68;
sine[36686]=-68;
sine[36687]=-68;
sine[36688]=-68;
sine[36689]=-68;
sine[36690]=-68;
sine[36691]=-68;
sine[36692]=-68;
sine[36693]=-68;
sine[36694]=-68;
sine[36695]=-68;
sine[36696]=-68;
sine[36697]=-68;
sine[36698]=-68;
sine[36699]=-68;
sine[36700]=-68;
sine[36701]=-68;
sine[36702]=-69;
sine[36703]=-69;
sine[36704]=-69;
sine[36705]=-69;
sine[36706]=-69;
sine[36707]=-69;
sine[36708]=-69;
sine[36709]=-69;
sine[36710]=-69;
sine[36711]=-69;
sine[36712]=-69;
sine[36713]=-69;
sine[36714]=-69;
sine[36715]=-69;
sine[36716]=-69;
sine[36717]=-69;
sine[36718]=-69;
sine[36719]=-69;
sine[36720]=-69;
sine[36721]=-69;
sine[36722]=-69;
sine[36723]=-69;
sine[36724]=-69;
sine[36725]=-69;
sine[36726]=-69;
sine[36727]=-69;
sine[36728]=-69;
sine[36729]=-69;
sine[36730]=-69;
sine[36731]=-69;
sine[36732]=-69;
sine[36733]=-69;
sine[36734]=-69;
sine[36735]=-69;
sine[36736]=-69;
sine[36737]=-69;
sine[36738]=-69;
sine[36739]=-69;
sine[36740]=-69;
sine[36741]=-69;
sine[36742]=-69;
sine[36743]=-69;
sine[36744]=-69;
sine[36745]=-69;
sine[36746]=-70;
sine[36747]=-70;
sine[36748]=-70;
sine[36749]=-70;
sine[36750]=-70;
sine[36751]=-70;
sine[36752]=-70;
sine[36753]=-70;
sine[36754]=-70;
sine[36755]=-70;
sine[36756]=-70;
sine[36757]=-70;
sine[36758]=-70;
sine[36759]=-70;
sine[36760]=-70;
sine[36761]=-70;
sine[36762]=-70;
sine[36763]=-70;
sine[36764]=-70;
sine[36765]=-70;
sine[36766]=-70;
sine[36767]=-70;
sine[36768]=-70;
sine[36769]=-70;
sine[36770]=-70;
sine[36771]=-70;
sine[36772]=-70;
sine[36773]=-70;
sine[36774]=-70;
sine[36775]=-70;
sine[36776]=-70;
sine[36777]=-70;
sine[36778]=-70;
sine[36779]=-70;
sine[36780]=-70;
sine[36781]=-70;
sine[36782]=-70;
sine[36783]=-70;
sine[36784]=-70;
sine[36785]=-70;
sine[36786]=-70;
sine[36787]=-70;
sine[36788]=-70;
sine[36789]=-70;
sine[36790]=-70;
sine[36791]=-71;
sine[36792]=-71;
sine[36793]=-71;
sine[36794]=-71;
sine[36795]=-71;
sine[36796]=-71;
sine[36797]=-71;
sine[36798]=-71;
sine[36799]=-71;
sine[36800]=-71;
sine[36801]=-71;
sine[36802]=-71;
sine[36803]=-71;
sine[36804]=-71;
sine[36805]=-71;
sine[36806]=-71;
sine[36807]=-71;
sine[36808]=-71;
sine[36809]=-71;
sine[36810]=-71;
sine[36811]=-71;
sine[36812]=-71;
sine[36813]=-71;
sine[36814]=-71;
sine[36815]=-71;
sine[36816]=-71;
sine[36817]=-71;
sine[36818]=-71;
sine[36819]=-71;
sine[36820]=-71;
sine[36821]=-71;
sine[36822]=-71;
sine[36823]=-71;
sine[36824]=-71;
sine[36825]=-71;
sine[36826]=-71;
sine[36827]=-71;
sine[36828]=-71;
sine[36829]=-71;
sine[36830]=-71;
sine[36831]=-71;
sine[36832]=-71;
sine[36833]=-71;
sine[36834]=-71;
sine[36835]=-71;
sine[36836]=-71;
sine[36837]=-71;
sine[36838]=-71;
sine[36839]=-71;
sine[36840]=-72;
sine[36841]=-72;
sine[36842]=-72;
sine[36843]=-72;
sine[36844]=-72;
sine[36845]=-72;
sine[36846]=-72;
sine[36847]=-72;
sine[36848]=-72;
sine[36849]=-72;
sine[36850]=-72;
sine[36851]=-72;
sine[36852]=-72;
sine[36853]=-72;
sine[36854]=-72;
sine[36855]=-72;
sine[36856]=-72;
sine[36857]=-72;
sine[36858]=-72;
sine[36859]=-72;
sine[36860]=-72;
sine[36861]=-72;
sine[36862]=-72;
sine[36863]=-72;
sine[36864]=-72;
sine[36865]=-72;
sine[36866]=-72;
sine[36867]=-72;
sine[36868]=-72;
sine[36869]=-72;
sine[36870]=-72;
sine[36871]=-72;
sine[36872]=-72;
sine[36873]=-72;
sine[36874]=-72;
sine[36875]=-72;
sine[36876]=-72;
sine[36877]=-72;
sine[36878]=-72;
sine[36879]=-72;
sine[36880]=-72;
sine[36881]=-72;
sine[36882]=-72;
sine[36883]=-72;
sine[36884]=-72;
sine[36885]=-72;
sine[36886]=-72;
sine[36887]=-72;
sine[36888]=-72;
sine[36889]=-72;
sine[36890]=-72;
sine[36891]=-72;
sine[36892]=-72;
sine[36893]=-73;
sine[36894]=-73;
sine[36895]=-73;
sine[36896]=-73;
sine[36897]=-73;
sine[36898]=-73;
sine[36899]=-73;
sine[36900]=-73;
sine[36901]=-73;
sine[36902]=-73;
sine[36903]=-73;
sine[36904]=-73;
sine[36905]=-73;
sine[36906]=-73;
sine[36907]=-73;
sine[36908]=-73;
sine[36909]=-73;
sine[36910]=-73;
sine[36911]=-73;
sine[36912]=-73;
sine[36913]=-73;
sine[36914]=-73;
sine[36915]=-73;
sine[36916]=-73;
sine[36917]=-73;
sine[36918]=-73;
sine[36919]=-73;
sine[36920]=-73;
sine[36921]=-73;
sine[36922]=-73;
sine[36923]=-73;
sine[36924]=-73;
sine[36925]=-73;
sine[36926]=-73;
sine[36927]=-73;
sine[36928]=-73;
sine[36929]=-73;
sine[36930]=-73;
sine[36931]=-73;
sine[36932]=-73;
sine[36933]=-73;
sine[36934]=-73;
sine[36935]=-73;
sine[36936]=-73;
sine[36937]=-73;
sine[36938]=-73;
sine[36939]=-73;
sine[36940]=-73;
sine[36941]=-73;
sine[36942]=-73;
sine[36943]=-73;
sine[36944]=-73;
sine[36945]=-73;
sine[36946]=-73;
sine[36947]=-73;
sine[36948]=-73;
sine[36949]=-73;
sine[36950]=-74;
sine[36951]=-74;
sine[36952]=-74;
sine[36953]=-74;
sine[36954]=-74;
sine[36955]=-74;
sine[36956]=-74;
sine[36957]=-74;
sine[36958]=-74;
sine[36959]=-74;
sine[36960]=-74;
sine[36961]=-74;
sine[36962]=-74;
sine[36963]=-74;
sine[36964]=-74;
sine[36965]=-74;
sine[36966]=-74;
sine[36967]=-74;
sine[36968]=-74;
sine[36969]=-74;
sine[36970]=-74;
sine[36971]=-74;
sine[36972]=-74;
sine[36973]=-74;
sine[36974]=-74;
sine[36975]=-74;
sine[36976]=-74;
sine[36977]=-74;
sine[36978]=-74;
sine[36979]=-74;
sine[36980]=-74;
sine[36981]=-74;
sine[36982]=-74;
sine[36983]=-74;
sine[36984]=-74;
sine[36985]=-74;
sine[36986]=-74;
sine[36987]=-74;
sine[36988]=-74;
sine[36989]=-74;
sine[36990]=-74;
sine[36991]=-74;
sine[36992]=-74;
sine[36993]=-74;
sine[36994]=-74;
sine[36995]=-74;
sine[36996]=-74;
sine[36997]=-74;
sine[36998]=-74;
sine[36999]=-74;
sine[37000]=-74;
sine[37001]=-74;
sine[37002]=-74;
sine[37003]=-74;
sine[37004]=-74;
sine[37005]=-74;
sine[37006]=-74;
sine[37007]=-74;
sine[37008]=-74;
sine[37009]=-74;
sine[37010]=-74;
sine[37011]=-74;
sine[37012]=-74;
sine[37013]=-74;
sine[37014]=-75;
sine[37015]=-75;
sine[37016]=-75;
sine[37017]=-75;
sine[37018]=-75;
sine[37019]=-75;
sine[37020]=-75;
sine[37021]=-75;
sine[37022]=-75;
sine[37023]=-75;
sine[37024]=-75;
sine[37025]=-75;
sine[37026]=-75;
sine[37027]=-75;
sine[37028]=-75;
sine[37029]=-75;
sine[37030]=-75;
sine[37031]=-75;
sine[37032]=-75;
sine[37033]=-75;
sine[37034]=-75;
sine[37035]=-75;
sine[37036]=-75;
sine[37037]=-75;
sine[37038]=-75;
sine[37039]=-75;
sine[37040]=-75;
sine[37041]=-75;
sine[37042]=-75;
sine[37043]=-75;
sine[37044]=-75;
sine[37045]=-75;
sine[37046]=-75;
sine[37047]=-75;
sine[37048]=-75;
sine[37049]=-75;
sine[37050]=-75;
sine[37051]=-75;
sine[37052]=-75;
sine[37053]=-75;
sine[37054]=-75;
sine[37055]=-75;
sine[37056]=-75;
sine[37057]=-75;
sine[37058]=-75;
sine[37059]=-75;
sine[37060]=-75;
sine[37061]=-75;
sine[37062]=-75;
sine[37063]=-75;
sine[37064]=-75;
sine[37065]=-75;
sine[37066]=-75;
sine[37067]=-75;
sine[37068]=-75;
sine[37069]=-75;
sine[37070]=-75;
sine[37071]=-75;
sine[37072]=-75;
sine[37073]=-75;
sine[37074]=-75;
sine[37075]=-75;
sine[37076]=-75;
sine[37077]=-75;
sine[37078]=-75;
sine[37079]=-75;
sine[37080]=-75;
sine[37081]=-75;
sine[37082]=-75;
sine[37083]=-75;
sine[37084]=-75;
sine[37085]=-75;
sine[37086]=-75;
sine[37087]=-76;
sine[37088]=-76;
sine[37089]=-76;
sine[37090]=-76;
sine[37091]=-76;
sine[37092]=-76;
sine[37093]=-76;
sine[37094]=-76;
sine[37095]=-76;
sine[37096]=-76;
sine[37097]=-76;
sine[37098]=-76;
sine[37099]=-76;
sine[37100]=-76;
sine[37101]=-76;
sine[37102]=-76;
sine[37103]=-76;
sine[37104]=-76;
sine[37105]=-76;
sine[37106]=-76;
sine[37107]=-76;
sine[37108]=-76;
sine[37109]=-76;
sine[37110]=-76;
sine[37111]=-76;
sine[37112]=-76;
sine[37113]=-76;
sine[37114]=-76;
sine[37115]=-76;
sine[37116]=-76;
sine[37117]=-76;
sine[37118]=-76;
sine[37119]=-76;
sine[37120]=-76;
sine[37121]=-76;
sine[37122]=-76;
sine[37123]=-76;
sine[37124]=-76;
sine[37125]=-76;
sine[37126]=-76;
sine[37127]=-76;
sine[37128]=-76;
sine[37129]=-76;
sine[37130]=-76;
sine[37131]=-76;
sine[37132]=-76;
sine[37133]=-76;
sine[37134]=-76;
sine[37135]=-76;
sine[37136]=-76;
sine[37137]=-76;
sine[37138]=-76;
sine[37139]=-76;
sine[37140]=-76;
sine[37141]=-76;
sine[37142]=-76;
sine[37143]=-76;
sine[37144]=-76;
sine[37145]=-76;
sine[37146]=-76;
sine[37147]=-76;
sine[37148]=-76;
sine[37149]=-76;
sine[37150]=-76;
sine[37151]=-76;
sine[37152]=-76;
sine[37153]=-76;
sine[37154]=-76;
sine[37155]=-76;
sine[37156]=-76;
sine[37157]=-76;
sine[37158]=-76;
sine[37159]=-76;
sine[37160]=-76;
sine[37161]=-76;
sine[37162]=-76;
sine[37163]=-76;
sine[37164]=-76;
sine[37165]=-76;
sine[37166]=-76;
sine[37167]=-76;
sine[37168]=-76;
sine[37169]=-76;
sine[37170]=-76;
sine[37171]=-76;
sine[37172]=-76;
sine[37173]=-76;
sine[37174]=-76;
sine[37175]=-77;
sine[37176]=-77;
sine[37177]=-77;
sine[37178]=-77;
sine[37179]=-77;
sine[37180]=-77;
sine[37181]=-77;
sine[37182]=-77;
sine[37183]=-77;
sine[37184]=-77;
sine[37185]=-77;
sine[37186]=-77;
sine[37187]=-77;
sine[37188]=-77;
sine[37189]=-77;
sine[37190]=-77;
sine[37191]=-77;
sine[37192]=-77;
sine[37193]=-77;
sine[37194]=-77;
sine[37195]=-77;
sine[37196]=-77;
sine[37197]=-77;
sine[37198]=-77;
sine[37199]=-77;
sine[37200]=-77;
sine[37201]=-77;
sine[37202]=-77;
sine[37203]=-77;
sine[37204]=-77;
sine[37205]=-77;
sine[37206]=-77;
sine[37207]=-77;
sine[37208]=-77;
sine[37209]=-77;
sine[37210]=-77;
sine[37211]=-77;
sine[37212]=-77;
sine[37213]=-77;
sine[37214]=-77;
sine[37215]=-77;
sine[37216]=-77;
sine[37217]=-77;
sine[37218]=-77;
sine[37219]=-77;
sine[37220]=-77;
sine[37221]=-77;
sine[37222]=-77;
sine[37223]=-77;
sine[37224]=-77;
sine[37225]=-77;
sine[37226]=-77;
sine[37227]=-77;
sine[37228]=-77;
sine[37229]=-77;
sine[37230]=-77;
sine[37231]=-77;
sine[37232]=-77;
sine[37233]=-77;
sine[37234]=-77;
sine[37235]=-77;
sine[37236]=-77;
sine[37237]=-77;
sine[37238]=-77;
sine[37239]=-77;
sine[37240]=-77;
sine[37241]=-77;
sine[37242]=-77;
sine[37243]=-77;
sine[37244]=-77;
sine[37245]=-77;
sine[37246]=-77;
sine[37247]=-77;
sine[37248]=-77;
sine[37249]=-77;
sine[37250]=-77;
sine[37251]=-77;
sine[37252]=-77;
sine[37253]=-77;
sine[37254]=-77;
sine[37255]=-77;
sine[37256]=-77;
sine[37257]=-77;
sine[37258]=-77;
sine[37259]=-77;
sine[37260]=-77;
sine[37261]=-77;
sine[37262]=-77;
sine[37263]=-77;
sine[37264]=-77;
sine[37265]=-77;
sine[37266]=-77;
sine[37267]=-77;
sine[37268]=-77;
sine[37269]=-77;
sine[37270]=-77;
sine[37271]=-77;
sine[37272]=-77;
sine[37273]=-77;
sine[37274]=-77;
sine[37275]=-77;
sine[37276]=-77;
sine[37277]=-77;
sine[37278]=-77;
sine[37279]=-77;
sine[37280]=-77;
sine[37281]=-77;
sine[37282]=-77;
sine[37283]=-77;
sine[37284]=-77;
sine[37285]=-77;
sine[37286]=-77;
sine[37287]=-77;
sine[37288]=-77;
sine[37289]=-77;
sine[37290]=-77;
sine[37291]=-77;
sine[37292]=-77;
sine[37293]=-77;
sine[37294]=-77;
sine[37295]=-77;
sine[37296]=-77;
sine[37297]=-77;
sine[37298]=-77;
sine[37299]=-78;
sine[37300]=-78;
sine[37301]=-78;
sine[37302]=-78;
sine[37303]=-78;
sine[37304]=-78;
sine[37305]=-78;
sine[37306]=-78;
sine[37307]=-78;
sine[37308]=-78;
sine[37309]=-78;
sine[37310]=-78;
sine[37311]=-78;
sine[37312]=-78;
sine[37313]=-78;
sine[37314]=-78;
sine[37315]=-78;
sine[37316]=-78;
sine[37317]=-78;
sine[37318]=-78;
sine[37319]=-78;
sine[37320]=-78;
sine[37321]=-78;
sine[37322]=-78;
sine[37323]=-78;
sine[37324]=-78;
sine[37325]=-78;
sine[37326]=-78;
sine[37327]=-78;
sine[37328]=-78;
sine[37329]=-78;
sine[37330]=-78;
sine[37331]=-78;
sine[37332]=-78;
sine[37333]=-78;
sine[37334]=-78;
sine[37335]=-78;
sine[37336]=-78;
sine[37337]=-78;
sine[37338]=-78;
sine[37339]=-78;
sine[37340]=-78;
sine[37341]=-78;
sine[37342]=-78;
sine[37343]=-78;
sine[37344]=-78;
sine[37345]=-78;
sine[37346]=-78;
sine[37347]=-78;
sine[37348]=-78;
sine[37349]=-78;
sine[37350]=-78;
sine[37351]=-78;
sine[37352]=-78;
sine[37353]=-78;
sine[37354]=-78;
sine[37355]=-78;
sine[37356]=-78;
sine[37357]=-78;
sine[37358]=-78;
sine[37359]=-78;
sine[37360]=-78;
sine[37361]=-78;
sine[37362]=-78;
sine[37363]=-78;
sine[37364]=-78;
sine[37365]=-78;
sine[37366]=-78;
sine[37367]=-78;
sine[37368]=-78;
sine[37369]=-78;
sine[37370]=-78;
sine[37371]=-78;
sine[37372]=-78;
sine[37373]=-78;
sine[37374]=-78;
sine[37375]=-78;
sine[37376]=-78;
sine[37377]=-78;
sine[37378]=-78;
sine[37379]=-78;
sine[37380]=-78;
sine[37381]=-78;
sine[37382]=-78;
sine[37383]=-78;
sine[37384]=-78;
sine[37385]=-78;
sine[37386]=-78;
sine[37387]=-78;
sine[37388]=-78;
sine[37389]=-78;
sine[37390]=-78;
sine[37391]=-78;
sine[37392]=-78;
sine[37393]=-78;
sine[37394]=-78;
sine[37395]=-78;
sine[37396]=-78;
sine[37397]=-78;
sine[37398]=-78;
sine[37399]=-78;
sine[37400]=-78;
sine[37401]=-78;
sine[37402]=-78;
sine[37403]=-78;
sine[37404]=-78;
sine[37405]=-78;
sine[37406]=-78;
sine[37407]=-78;
sine[37408]=-78;
sine[37409]=-78;
sine[37410]=-78;
sine[37411]=-78;
sine[37412]=-78;
sine[37413]=-78;
sine[37414]=-78;
sine[37415]=-78;
sine[37416]=-78;
sine[37417]=-78;
sine[37418]=-78;
sine[37419]=-78;
sine[37420]=-78;
sine[37421]=-78;
sine[37422]=-78;
sine[37423]=-78;
sine[37424]=-78;
sine[37425]=-78;
sine[37426]=-78;
sine[37427]=-78;
sine[37428]=-78;
sine[37429]=-78;
sine[37430]=-78;
sine[37431]=-78;
sine[37432]=-78;
sine[37433]=-78;
sine[37434]=-78;
sine[37435]=-78;
sine[37436]=-78;
sine[37437]=-78;
sine[37438]=-78;
sine[37439]=-78;
sine[37440]=-78;
sine[37441]=-78;
sine[37442]=-78;
sine[37443]=-78;
sine[37444]=-78;
sine[37445]=-78;
sine[37446]=-78;
sine[37447]=-78;
sine[37448]=-78;
sine[37449]=-78;
sine[37450]=-78;
sine[37451]=-78;
sine[37452]=-78;
sine[37453]=-78;
sine[37454]=-78;
sine[37455]=-78;
sine[37456]=-78;
sine[37457]=-78;
sine[37458]=-78;
sine[37459]=-78;
sine[37460]=-78;
sine[37461]=-78;
sine[37462]=-78;
sine[37463]=-78;
sine[37464]=-78;
sine[37465]=-78;
sine[37466]=-78;
sine[37467]=-78;
sine[37468]=-78;
sine[37469]=-78;
sine[37470]=-78;
sine[37471]=-78;
sine[37472]=-78;
sine[37473]=-78;
sine[37474]=-78;
sine[37475]=-78;
sine[37476]=-78;
sine[37477]=-78;
sine[37478]=-78;
sine[37479]=-78;
sine[37480]=-78;
sine[37481]=-78;
sine[37482]=-78;
sine[37483]=-78;
sine[37484]=-78;
sine[37485]=-78;
sine[37486]=-78;
sine[37487]=-78;
sine[37488]=-78;
sine[37489]=-78;
sine[37490]=-78;
sine[37491]=-78;
sine[37492]=-78;
sine[37493]=-78;
sine[37494]=-78;
sine[37495]=-78;
sine[37496]=-78;
sine[37497]=-78;
sine[37498]=-78;
sine[37499]=-78;
sine[37500]=-78;
sine[37501]=-78;
sine[37502]=-78;
sine[37503]=-78;
sine[37504]=-78;
sine[37505]=-78;
sine[37506]=-78;
sine[37507]=-78;
sine[37508]=-78;
sine[37509]=-78;
sine[37510]=-78;
sine[37511]=-78;
sine[37512]=-78;
sine[37513]=-78;
sine[37514]=-78;
sine[37515]=-78;
sine[37516]=-78;
sine[37517]=-78;
sine[37518]=-78;
sine[37519]=-78;
sine[37520]=-78;
sine[37521]=-78;
sine[37522]=-78;
sine[37523]=-78;
sine[37524]=-78;
sine[37525]=-78;
sine[37526]=-78;
sine[37527]=-78;
sine[37528]=-78;
sine[37529]=-78;
sine[37530]=-78;
sine[37531]=-78;
sine[37532]=-78;
sine[37533]=-78;
sine[37534]=-78;
sine[37535]=-78;
sine[37536]=-78;
sine[37537]=-78;
sine[37538]=-78;
sine[37539]=-78;
sine[37540]=-78;
sine[37541]=-78;
sine[37542]=-78;
sine[37543]=-78;
sine[37544]=-78;
sine[37545]=-78;
sine[37546]=-78;
sine[37547]=-78;
sine[37548]=-78;
sine[37549]=-78;
sine[37550]=-78;
sine[37551]=-78;
sine[37552]=-78;
sine[37553]=-78;
sine[37554]=-78;
sine[37555]=-78;
sine[37556]=-78;
sine[37557]=-78;
sine[37558]=-78;
sine[37559]=-78;
sine[37560]=-78;
sine[37561]=-78;
sine[37562]=-78;
sine[37563]=-78;
sine[37564]=-78;
sine[37565]=-78;
sine[37566]=-78;
sine[37567]=-78;
sine[37568]=-78;
sine[37569]=-78;
sine[37570]=-78;
sine[37571]=-78;
sine[37572]=-78;
sine[37573]=-78;
sine[37574]=-78;
sine[37575]=-78;
sine[37576]=-78;
sine[37577]=-78;
sine[37578]=-78;
sine[37579]=-78;
sine[37580]=-78;
sine[37581]=-78;
sine[37582]=-78;
sine[37583]=-78;
sine[37584]=-78;
sine[37585]=-78;
sine[37586]=-78;
sine[37587]=-78;
sine[37588]=-78;
sine[37589]=-78;
sine[37590]=-78;
sine[37591]=-78;
sine[37592]=-78;
sine[37593]=-78;
sine[37594]=-78;
sine[37595]=-78;
sine[37596]=-78;
sine[37597]=-78;
sine[37598]=-78;
sine[37599]=-78;
sine[37600]=-78;
sine[37601]=-78;
sine[37602]=-78;
sine[37603]=-78;
sine[37604]=-78;
sine[37605]=-78;
sine[37606]=-78;
sine[37607]=-78;
sine[37608]=-78;
sine[37609]=-78;
sine[37610]=-78;
sine[37611]=-78;
sine[37612]=-78;
sine[37613]=-78;
sine[37614]=-78;
sine[37615]=-78;
sine[37616]=-78;
sine[37617]=-78;
sine[37618]=-78;
sine[37619]=-78;
sine[37620]=-78;
sine[37621]=-78;
sine[37622]=-78;
sine[37623]=-78;
sine[37624]=-78;
sine[37625]=-78;
sine[37626]=-78;
sine[37627]=-78;
sine[37628]=-78;
sine[37629]=-78;
sine[37630]=-78;
sine[37631]=-78;
sine[37632]=-78;
sine[37633]=-78;
sine[37634]=-78;
sine[37635]=-78;
sine[37636]=-78;
sine[37637]=-78;
sine[37638]=-78;
sine[37639]=-78;
sine[37640]=-78;
sine[37641]=-78;
sine[37642]=-78;
sine[37643]=-78;
sine[37644]=-78;
sine[37645]=-78;
sine[37646]=-78;
sine[37647]=-78;
sine[37648]=-78;
sine[37649]=-78;
sine[37650]=-78;
sine[37651]=-78;
sine[37652]=-78;
sine[37653]=-78;
sine[37654]=-78;
sine[37655]=-78;
sine[37656]=-78;
sine[37657]=-78;
sine[37658]=-78;
sine[37659]=-78;
sine[37660]=-78;
sine[37661]=-78;
sine[37662]=-78;
sine[37663]=-78;
sine[37664]=-78;
sine[37665]=-78;
sine[37666]=-78;
sine[37667]=-78;
sine[37668]=-78;
sine[37669]=-78;
sine[37670]=-78;
sine[37671]=-78;
sine[37672]=-78;
sine[37673]=-78;
sine[37674]=-78;
sine[37675]=-78;
sine[37676]=-78;
sine[37677]=-78;
sine[37678]=-78;
sine[37679]=-78;
sine[37680]=-78;
sine[37681]=-78;
sine[37682]=-78;
sine[37683]=-78;
sine[37684]=-78;
sine[37685]=-78;
sine[37686]=-78;
sine[37687]=-78;
sine[37688]=-78;
sine[37689]=-78;
sine[37690]=-78;
sine[37691]=-78;
sine[37692]=-78;
sine[37693]=-78;
sine[37694]=-78;
sine[37695]=-78;
sine[37696]=-78;
sine[37697]=-78;
sine[37698]=-78;
sine[37699]=-78;
sine[37700]=-78;
sine[37701]=-78;
sine[37702]=-77;
sine[37703]=-77;
sine[37704]=-77;
sine[37705]=-77;
sine[37706]=-77;
sine[37707]=-77;
sine[37708]=-77;
sine[37709]=-77;
sine[37710]=-77;
sine[37711]=-77;
sine[37712]=-77;
sine[37713]=-77;
sine[37714]=-77;
sine[37715]=-77;
sine[37716]=-77;
sine[37717]=-77;
sine[37718]=-77;
sine[37719]=-77;
sine[37720]=-77;
sine[37721]=-77;
sine[37722]=-77;
sine[37723]=-77;
sine[37724]=-77;
sine[37725]=-77;
sine[37726]=-77;
sine[37727]=-77;
sine[37728]=-77;
sine[37729]=-77;
sine[37730]=-77;
sine[37731]=-77;
sine[37732]=-77;
sine[37733]=-77;
sine[37734]=-77;
sine[37735]=-77;
sine[37736]=-77;
sine[37737]=-77;
sine[37738]=-77;
sine[37739]=-77;
sine[37740]=-77;
sine[37741]=-77;
sine[37742]=-77;
sine[37743]=-77;
sine[37744]=-77;
sine[37745]=-77;
sine[37746]=-77;
sine[37747]=-77;
sine[37748]=-77;
sine[37749]=-77;
sine[37750]=-77;
sine[37751]=-77;
sine[37752]=-77;
sine[37753]=-77;
sine[37754]=-77;
sine[37755]=-77;
sine[37756]=-77;
sine[37757]=-77;
sine[37758]=-77;
sine[37759]=-77;
sine[37760]=-77;
sine[37761]=-77;
sine[37762]=-77;
sine[37763]=-77;
sine[37764]=-77;
sine[37765]=-77;
sine[37766]=-77;
sine[37767]=-77;
sine[37768]=-77;
sine[37769]=-77;
sine[37770]=-77;
sine[37771]=-77;
sine[37772]=-77;
sine[37773]=-77;
sine[37774]=-77;
sine[37775]=-77;
sine[37776]=-77;
sine[37777]=-77;
sine[37778]=-77;
sine[37779]=-77;
sine[37780]=-77;
sine[37781]=-77;
sine[37782]=-77;
sine[37783]=-77;
sine[37784]=-77;
sine[37785]=-77;
sine[37786]=-77;
sine[37787]=-77;
sine[37788]=-77;
sine[37789]=-77;
sine[37790]=-77;
sine[37791]=-77;
sine[37792]=-77;
sine[37793]=-77;
sine[37794]=-77;
sine[37795]=-77;
sine[37796]=-77;
sine[37797]=-77;
sine[37798]=-77;
sine[37799]=-77;
sine[37800]=-77;
sine[37801]=-77;
sine[37802]=-77;
sine[37803]=-77;
sine[37804]=-77;
sine[37805]=-77;
sine[37806]=-77;
sine[37807]=-77;
sine[37808]=-77;
sine[37809]=-77;
sine[37810]=-77;
sine[37811]=-77;
sine[37812]=-77;
sine[37813]=-77;
sine[37814]=-77;
sine[37815]=-77;
sine[37816]=-77;
sine[37817]=-77;
sine[37818]=-77;
sine[37819]=-77;
sine[37820]=-77;
sine[37821]=-77;
sine[37822]=-77;
sine[37823]=-77;
sine[37824]=-77;
sine[37825]=-77;
sine[37826]=-76;
sine[37827]=-76;
sine[37828]=-76;
sine[37829]=-76;
sine[37830]=-76;
sine[37831]=-76;
sine[37832]=-76;
sine[37833]=-76;
sine[37834]=-76;
sine[37835]=-76;
sine[37836]=-76;
sine[37837]=-76;
sine[37838]=-76;
sine[37839]=-76;
sine[37840]=-76;
sine[37841]=-76;
sine[37842]=-76;
sine[37843]=-76;
sine[37844]=-76;
sine[37845]=-76;
sine[37846]=-76;
sine[37847]=-76;
sine[37848]=-76;
sine[37849]=-76;
sine[37850]=-76;
sine[37851]=-76;
sine[37852]=-76;
sine[37853]=-76;
sine[37854]=-76;
sine[37855]=-76;
sine[37856]=-76;
sine[37857]=-76;
sine[37858]=-76;
sine[37859]=-76;
sine[37860]=-76;
sine[37861]=-76;
sine[37862]=-76;
sine[37863]=-76;
sine[37864]=-76;
sine[37865]=-76;
sine[37866]=-76;
sine[37867]=-76;
sine[37868]=-76;
sine[37869]=-76;
sine[37870]=-76;
sine[37871]=-76;
sine[37872]=-76;
sine[37873]=-76;
sine[37874]=-76;
sine[37875]=-76;
sine[37876]=-76;
sine[37877]=-76;
sine[37878]=-76;
sine[37879]=-76;
sine[37880]=-76;
sine[37881]=-76;
sine[37882]=-76;
sine[37883]=-76;
sine[37884]=-76;
sine[37885]=-76;
sine[37886]=-76;
sine[37887]=-76;
sine[37888]=-76;
sine[37889]=-76;
sine[37890]=-76;
sine[37891]=-76;
sine[37892]=-76;
sine[37893]=-76;
sine[37894]=-76;
sine[37895]=-76;
sine[37896]=-76;
sine[37897]=-76;
sine[37898]=-76;
sine[37899]=-76;
sine[37900]=-76;
sine[37901]=-76;
sine[37902]=-76;
sine[37903]=-76;
sine[37904]=-76;
sine[37905]=-76;
sine[37906]=-76;
sine[37907]=-76;
sine[37908]=-76;
sine[37909]=-76;
sine[37910]=-76;
sine[37911]=-76;
sine[37912]=-76;
sine[37913]=-76;
sine[37914]=-75;
sine[37915]=-75;
sine[37916]=-75;
sine[37917]=-75;
sine[37918]=-75;
sine[37919]=-75;
sine[37920]=-75;
sine[37921]=-75;
sine[37922]=-75;
sine[37923]=-75;
sine[37924]=-75;
sine[37925]=-75;
sine[37926]=-75;
sine[37927]=-75;
sine[37928]=-75;
sine[37929]=-75;
sine[37930]=-75;
sine[37931]=-75;
sine[37932]=-75;
sine[37933]=-75;
sine[37934]=-75;
sine[37935]=-75;
sine[37936]=-75;
sine[37937]=-75;
sine[37938]=-75;
sine[37939]=-75;
sine[37940]=-75;
sine[37941]=-75;
sine[37942]=-75;
sine[37943]=-75;
sine[37944]=-75;
sine[37945]=-75;
sine[37946]=-75;
sine[37947]=-75;
sine[37948]=-75;
sine[37949]=-75;
sine[37950]=-75;
sine[37951]=-75;
sine[37952]=-75;
sine[37953]=-75;
sine[37954]=-75;
sine[37955]=-75;
sine[37956]=-75;
sine[37957]=-75;
sine[37958]=-75;
sine[37959]=-75;
sine[37960]=-75;
sine[37961]=-75;
sine[37962]=-75;
sine[37963]=-75;
sine[37964]=-75;
sine[37965]=-75;
sine[37966]=-75;
sine[37967]=-75;
sine[37968]=-75;
sine[37969]=-75;
sine[37970]=-75;
sine[37971]=-75;
sine[37972]=-75;
sine[37973]=-75;
sine[37974]=-75;
sine[37975]=-75;
sine[37976]=-75;
sine[37977]=-75;
sine[37978]=-75;
sine[37979]=-75;
sine[37980]=-75;
sine[37981]=-75;
sine[37982]=-75;
sine[37983]=-75;
sine[37984]=-75;
sine[37985]=-75;
sine[37986]=-75;
sine[37987]=-74;
sine[37988]=-74;
sine[37989]=-74;
sine[37990]=-74;
sine[37991]=-74;
sine[37992]=-74;
sine[37993]=-74;
sine[37994]=-74;
sine[37995]=-74;
sine[37996]=-74;
sine[37997]=-74;
sine[37998]=-74;
sine[37999]=-74;
sine[38000]=-74;
sine[38001]=-74;
sine[38002]=-74;
sine[38003]=-74;
sine[38004]=-74;
sine[38005]=-74;
sine[38006]=-74;
sine[38007]=-74;
sine[38008]=-74;
sine[38009]=-74;
sine[38010]=-74;
sine[38011]=-74;
sine[38012]=-74;
sine[38013]=-74;
sine[38014]=-74;
sine[38015]=-74;
sine[38016]=-74;
sine[38017]=-74;
sine[38018]=-74;
sine[38019]=-74;
sine[38020]=-74;
sine[38021]=-74;
sine[38022]=-74;
sine[38023]=-74;
sine[38024]=-74;
sine[38025]=-74;
sine[38026]=-74;
sine[38027]=-74;
sine[38028]=-74;
sine[38029]=-74;
sine[38030]=-74;
sine[38031]=-74;
sine[38032]=-74;
sine[38033]=-74;
sine[38034]=-74;
sine[38035]=-74;
sine[38036]=-74;
sine[38037]=-74;
sine[38038]=-74;
sine[38039]=-74;
sine[38040]=-74;
sine[38041]=-74;
sine[38042]=-74;
sine[38043]=-74;
sine[38044]=-74;
sine[38045]=-74;
sine[38046]=-74;
sine[38047]=-74;
sine[38048]=-74;
sine[38049]=-74;
sine[38050]=-74;
sine[38051]=-73;
sine[38052]=-73;
sine[38053]=-73;
sine[38054]=-73;
sine[38055]=-73;
sine[38056]=-73;
sine[38057]=-73;
sine[38058]=-73;
sine[38059]=-73;
sine[38060]=-73;
sine[38061]=-73;
sine[38062]=-73;
sine[38063]=-73;
sine[38064]=-73;
sine[38065]=-73;
sine[38066]=-73;
sine[38067]=-73;
sine[38068]=-73;
sine[38069]=-73;
sine[38070]=-73;
sine[38071]=-73;
sine[38072]=-73;
sine[38073]=-73;
sine[38074]=-73;
sine[38075]=-73;
sine[38076]=-73;
sine[38077]=-73;
sine[38078]=-73;
sine[38079]=-73;
sine[38080]=-73;
sine[38081]=-73;
sine[38082]=-73;
sine[38083]=-73;
sine[38084]=-73;
sine[38085]=-73;
sine[38086]=-73;
sine[38087]=-73;
sine[38088]=-73;
sine[38089]=-73;
sine[38090]=-73;
sine[38091]=-73;
sine[38092]=-73;
sine[38093]=-73;
sine[38094]=-73;
sine[38095]=-73;
sine[38096]=-73;
sine[38097]=-73;
sine[38098]=-73;
sine[38099]=-73;
sine[38100]=-73;
sine[38101]=-73;
sine[38102]=-73;
sine[38103]=-73;
sine[38104]=-73;
sine[38105]=-73;
sine[38106]=-73;
sine[38107]=-73;
sine[38108]=-72;
sine[38109]=-72;
sine[38110]=-72;
sine[38111]=-72;
sine[38112]=-72;
sine[38113]=-72;
sine[38114]=-72;
sine[38115]=-72;
sine[38116]=-72;
sine[38117]=-72;
sine[38118]=-72;
sine[38119]=-72;
sine[38120]=-72;
sine[38121]=-72;
sine[38122]=-72;
sine[38123]=-72;
sine[38124]=-72;
sine[38125]=-72;
sine[38126]=-72;
sine[38127]=-72;
sine[38128]=-72;
sine[38129]=-72;
sine[38130]=-72;
sine[38131]=-72;
sine[38132]=-72;
sine[38133]=-72;
sine[38134]=-72;
sine[38135]=-72;
sine[38136]=-72;
sine[38137]=-72;
sine[38138]=-72;
sine[38139]=-72;
sine[38140]=-72;
sine[38141]=-72;
sine[38142]=-72;
sine[38143]=-72;
sine[38144]=-72;
sine[38145]=-72;
sine[38146]=-72;
sine[38147]=-72;
sine[38148]=-72;
sine[38149]=-72;
sine[38150]=-72;
sine[38151]=-72;
sine[38152]=-72;
sine[38153]=-72;
sine[38154]=-72;
sine[38155]=-72;
sine[38156]=-72;
sine[38157]=-72;
sine[38158]=-72;
sine[38159]=-72;
sine[38160]=-72;
sine[38161]=-71;
sine[38162]=-71;
sine[38163]=-71;
sine[38164]=-71;
sine[38165]=-71;
sine[38166]=-71;
sine[38167]=-71;
sine[38168]=-71;
sine[38169]=-71;
sine[38170]=-71;
sine[38171]=-71;
sine[38172]=-71;
sine[38173]=-71;
sine[38174]=-71;
sine[38175]=-71;
sine[38176]=-71;
sine[38177]=-71;
sine[38178]=-71;
sine[38179]=-71;
sine[38180]=-71;
sine[38181]=-71;
sine[38182]=-71;
sine[38183]=-71;
sine[38184]=-71;
sine[38185]=-71;
sine[38186]=-71;
sine[38187]=-71;
sine[38188]=-71;
sine[38189]=-71;
sine[38190]=-71;
sine[38191]=-71;
sine[38192]=-71;
sine[38193]=-71;
sine[38194]=-71;
sine[38195]=-71;
sine[38196]=-71;
sine[38197]=-71;
sine[38198]=-71;
sine[38199]=-71;
sine[38200]=-71;
sine[38201]=-71;
sine[38202]=-71;
sine[38203]=-71;
sine[38204]=-71;
sine[38205]=-71;
sine[38206]=-71;
sine[38207]=-71;
sine[38208]=-71;
sine[38209]=-71;
sine[38210]=-70;
sine[38211]=-70;
sine[38212]=-70;
sine[38213]=-70;
sine[38214]=-70;
sine[38215]=-70;
sine[38216]=-70;
sine[38217]=-70;
sine[38218]=-70;
sine[38219]=-70;
sine[38220]=-70;
sine[38221]=-70;
sine[38222]=-70;
sine[38223]=-70;
sine[38224]=-70;
sine[38225]=-70;
sine[38226]=-70;
sine[38227]=-70;
sine[38228]=-70;
sine[38229]=-70;
sine[38230]=-70;
sine[38231]=-70;
sine[38232]=-70;
sine[38233]=-70;
sine[38234]=-70;
sine[38235]=-70;
sine[38236]=-70;
sine[38237]=-70;
sine[38238]=-70;
sine[38239]=-70;
sine[38240]=-70;
sine[38241]=-70;
sine[38242]=-70;
sine[38243]=-70;
sine[38244]=-70;
sine[38245]=-70;
sine[38246]=-70;
sine[38247]=-70;
sine[38248]=-70;
sine[38249]=-70;
sine[38250]=-70;
sine[38251]=-70;
sine[38252]=-70;
sine[38253]=-70;
sine[38254]=-70;
sine[38255]=-69;
sine[38256]=-69;
sine[38257]=-69;
sine[38258]=-69;
sine[38259]=-69;
sine[38260]=-69;
sine[38261]=-69;
sine[38262]=-69;
sine[38263]=-69;
sine[38264]=-69;
sine[38265]=-69;
sine[38266]=-69;
sine[38267]=-69;
sine[38268]=-69;
sine[38269]=-69;
sine[38270]=-69;
sine[38271]=-69;
sine[38272]=-69;
sine[38273]=-69;
sine[38274]=-69;
sine[38275]=-69;
sine[38276]=-69;
sine[38277]=-69;
sine[38278]=-69;
sine[38279]=-69;
sine[38280]=-69;
sine[38281]=-69;
sine[38282]=-69;
sine[38283]=-69;
sine[38284]=-69;
sine[38285]=-69;
sine[38286]=-69;
sine[38287]=-69;
sine[38288]=-69;
sine[38289]=-69;
sine[38290]=-69;
sine[38291]=-69;
sine[38292]=-69;
sine[38293]=-69;
sine[38294]=-69;
sine[38295]=-69;
sine[38296]=-69;
sine[38297]=-69;
sine[38298]=-69;
sine[38299]=-68;
sine[38300]=-68;
sine[38301]=-68;
sine[38302]=-68;
sine[38303]=-68;
sine[38304]=-68;
sine[38305]=-68;
sine[38306]=-68;
sine[38307]=-68;
sine[38308]=-68;
sine[38309]=-68;
sine[38310]=-68;
sine[38311]=-68;
sine[38312]=-68;
sine[38313]=-68;
sine[38314]=-68;
sine[38315]=-68;
sine[38316]=-68;
sine[38317]=-68;
sine[38318]=-68;
sine[38319]=-68;
sine[38320]=-68;
sine[38321]=-68;
sine[38322]=-68;
sine[38323]=-68;
sine[38324]=-68;
sine[38325]=-68;
sine[38326]=-68;
sine[38327]=-68;
sine[38328]=-68;
sine[38329]=-68;
sine[38330]=-68;
sine[38331]=-68;
sine[38332]=-68;
sine[38333]=-68;
sine[38334]=-68;
sine[38335]=-68;
sine[38336]=-68;
sine[38337]=-68;
sine[38338]=-68;
sine[38339]=-68;
sine[38340]=-67;
sine[38341]=-67;
sine[38342]=-67;
sine[38343]=-67;
sine[38344]=-67;
sine[38345]=-67;
sine[38346]=-67;
sine[38347]=-67;
sine[38348]=-67;
sine[38349]=-67;
sine[38350]=-67;
sine[38351]=-67;
sine[38352]=-67;
sine[38353]=-67;
sine[38354]=-67;
sine[38355]=-67;
sine[38356]=-67;
sine[38357]=-67;
sine[38358]=-67;
sine[38359]=-67;
sine[38360]=-67;
sine[38361]=-67;
sine[38362]=-67;
sine[38363]=-67;
sine[38364]=-67;
sine[38365]=-67;
sine[38366]=-67;
sine[38367]=-67;
sine[38368]=-67;
sine[38369]=-67;
sine[38370]=-67;
sine[38371]=-67;
sine[38372]=-67;
sine[38373]=-67;
sine[38374]=-67;
sine[38375]=-67;
sine[38376]=-67;
sine[38377]=-67;
sine[38378]=-67;
sine[38379]=-67;
sine[38380]=-66;
sine[38381]=-66;
sine[38382]=-66;
sine[38383]=-66;
sine[38384]=-66;
sine[38385]=-66;
sine[38386]=-66;
sine[38387]=-66;
sine[38388]=-66;
sine[38389]=-66;
sine[38390]=-66;
sine[38391]=-66;
sine[38392]=-66;
sine[38393]=-66;
sine[38394]=-66;
sine[38395]=-66;
sine[38396]=-66;
sine[38397]=-66;
sine[38398]=-66;
sine[38399]=-66;
sine[38400]=-66;
sine[38401]=-66;
sine[38402]=-66;
sine[38403]=-66;
sine[38404]=-66;
sine[38405]=-66;
sine[38406]=-66;
sine[38407]=-66;
sine[38408]=-66;
sine[38409]=-66;
sine[38410]=-66;
sine[38411]=-66;
sine[38412]=-66;
sine[38413]=-66;
sine[38414]=-66;
sine[38415]=-66;
sine[38416]=-66;
sine[38417]=-66;
sine[38418]=-65;
sine[38419]=-65;
sine[38420]=-65;
sine[38421]=-65;
sine[38422]=-65;
sine[38423]=-65;
sine[38424]=-65;
sine[38425]=-65;
sine[38426]=-65;
sine[38427]=-65;
sine[38428]=-65;
sine[38429]=-65;
sine[38430]=-65;
sine[38431]=-65;
sine[38432]=-65;
sine[38433]=-65;
sine[38434]=-65;
sine[38435]=-65;
sine[38436]=-65;
sine[38437]=-65;
sine[38438]=-65;
sine[38439]=-65;
sine[38440]=-65;
sine[38441]=-65;
sine[38442]=-65;
sine[38443]=-65;
sine[38444]=-65;
sine[38445]=-65;
sine[38446]=-65;
sine[38447]=-65;
sine[38448]=-65;
sine[38449]=-65;
sine[38450]=-65;
sine[38451]=-65;
sine[38452]=-65;
sine[38453]=-65;
sine[38454]=-65;
sine[38455]=-64;
sine[38456]=-64;
sine[38457]=-64;
sine[38458]=-64;
sine[38459]=-64;
sine[38460]=-64;
sine[38461]=-64;
sine[38462]=-64;
sine[38463]=-64;
sine[38464]=-64;
sine[38465]=-64;
sine[38466]=-64;
sine[38467]=-64;
sine[38468]=-64;
sine[38469]=-64;
sine[38470]=-64;
sine[38471]=-64;
sine[38472]=-64;
sine[38473]=-64;
sine[38474]=-64;
sine[38475]=-64;
sine[38476]=-64;
sine[38477]=-64;
sine[38478]=-64;
sine[38479]=-64;
sine[38480]=-64;
sine[38481]=-64;
sine[38482]=-64;
sine[38483]=-64;
sine[38484]=-64;
sine[38485]=-64;
sine[38486]=-64;
sine[38487]=-64;
sine[38488]=-64;
sine[38489]=-64;
sine[38490]=-63;
sine[38491]=-63;
sine[38492]=-63;
sine[38493]=-63;
sine[38494]=-63;
sine[38495]=-63;
sine[38496]=-63;
sine[38497]=-63;
sine[38498]=-63;
sine[38499]=-63;
sine[38500]=-63;
sine[38501]=-63;
sine[38502]=-63;
sine[38503]=-63;
sine[38504]=-63;
sine[38505]=-63;
sine[38506]=-63;
sine[38507]=-63;
sine[38508]=-63;
sine[38509]=-63;
sine[38510]=-63;
sine[38511]=-63;
sine[38512]=-63;
sine[38513]=-63;
sine[38514]=-63;
sine[38515]=-63;
sine[38516]=-63;
sine[38517]=-63;
sine[38518]=-63;
sine[38519]=-63;
sine[38520]=-63;
sine[38521]=-63;
sine[38522]=-63;
sine[38523]=-63;
sine[38524]=-63;
sine[38525]=-62;
sine[38526]=-62;
sine[38527]=-62;
sine[38528]=-62;
sine[38529]=-62;
sine[38530]=-62;
sine[38531]=-62;
sine[38532]=-62;
sine[38533]=-62;
sine[38534]=-62;
sine[38535]=-62;
sine[38536]=-62;
sine[38537]=-62;
sine[38538]=-62;
sine[38539]=-62;
sine[38540]=-62;
sine[38541]=-62;
sine[38542]=-62;
sine[38543]=-62;
sine[38544]=-62;
sine[38545]=-62;
sine[38546]=-62;
sine[38547]=-62;
sine[38548]=-62;
sine[38549]=-62;
sine[38550]=-62;
sine[38551]=-62;
sine[38552]=-62;
sine[38553]=-62;
sine[38554]=-62;
sine[38555]=-62;
sine[38556]=-62;
sine[38557]=-62;
sine[38558]=-61;
sine[38559]=-61;
sine[38560]=-61;
sine[38561]=-61;
sine[38562]=-61;
sine[38563]=-61;
sine[38564]=-61;
sine[38565]=-61;
sine[38566]=-61;
sine[38567]=-61;
sine[38568]=-61;
sine[38569]=-61;
sine[38570]=-61;
sine[38571]=-61;
sine[38572]=-61;
sine[38573]=-61;
sine[38574]=-61;
sine[38575]=-61;
sine[38576]=-61;
sine[38577]=-61;
sine[38578]=-61;
sine[38579]=-61;
sine[38580]=-61;
sine[38581]=-61;
sine[38582]=-61;
sine[38583]=-61;
sine[38584]=-61;
sine[38585]=-61;
sine[38586]=-61;
sine[38587]=-61;
sine[38588]=-61;
sine[38589]=-61;
sine[38590]=-61;
sine[38591]=-60;
sine[38592]=-60;
sine[38593]=-60;
sine[38594]=-60;
sine[38595]=-60;
sine[38596]=-60;
sine[38597]=-60;
sine[38598]=-60;
sine[38599]=-60;
sine[38600]=-60;
sine[38601]=-60;
sine[38602]=-60;
sine[38603]=-60;
sine[38604]=-60;
sine[38605]=-60;
sine[38606]=-60;
sine[38607]=-60;
sine[38608]=-60;
sine[38609]=-60;
sine[38610]=-60;
sine[38611]=-60;
sine[38612]=-60;
sine[38613]=-60;
sine[38614]=-60;
sine[38615]=-60;
sine[38616]=-60;
sine[38617]=-60;
sine[38618]=-60;
sine[38619]=-60;
sine[38620]=-60;
sine[38621]=-60;
sine[38622]=-60;
sine[38623]=-59;
sine[38624]=-59;
sine[38625]=-59;
sine[38626]=-59;
sine[38627]=-59;
sine[38628]=-59;
sine[38629]=-59;
sine[38630]=-59;
sine[38631]=-59;
sine[38632]=-59;
sine[38633]=-59;
sine[38634]=-59;
sine[38635]=-59;
sine[38636]=-59;
sine[38637]=-59;
sine[38638]=-59;
sine[38639]=-59;
sine[38640]=-59;
sine[38641]=-59;
sine[38642]=-59;
sine[38643]=-59;
sine[38644]=-59;
sine[38645]=-59;
sine[38646]=-59;
sine[38647]=-59;
sine[38648]=-59;
sine[38649]=-59;
sine[38650]=-59;
sine[38651]=-59;
sine[38652]=-59;
sine[38653]=-59;
sine[38654]=-58;
sine[38655]=-58;
sine[38656]=-58;
sine[38657]=-58;
sine[38658]=-58;
sine[38659]=-58;
sine[38660]=-58;
sine[38661]=-58;
sine[38662]=-58;
sine[38663]=-58;
sine[38664]=-58;
sine[38665]=-58;
sine[38666]=-58;
sine[38667]=-58;
sine[38668]=-58;
sine[38669]=-58;
sine[38670]=-58;
sine[38671]=-58;
sine[38672]=-58;
sine[38673]=-58;
sine[38674]=-58;
sine[38675]=-58;
sine[38676]=-58;
sine[38677]=-58;
sine[38678]=-58;
sine[38679]=-58;
sine[38680]=-58;
sine[38681]=-58;
sine[38682]=-58;
sine[38683]=-58;
sine[38684]=-57;
sine[38685]=-57;
sine[38686]=-57;
sine[38687]=-57;
sine[38688]=-57;
sine[38689]=-57;
sine[38690]=-57;
sine[38691]=-57;
sine[38692]=-57;
sine[38693]=-57;
sine[38694]=-57;
sine[38695]=-57;
sine[38696]=-57;
sine[38697]=-57;
sine[38698]=-57;
sine[38699]=-57;
sine[38700]=-57;
sine[38701]=-57;
sine[38702]=-57;
sine[38703]=-57;
sine[38704]=-57;
sine[38705]=-57;
sine[38706]=-57;
sine[38707]=-57;
sine[38708]=-57;
sine[38709]=-57;
sine[38710]=-57;
sine[38711]=-57;
sine[38712]=-57;
sine[38713]=-57;
sine[38714]=-56;
sine[38715]=-56;
sine[38716]=-56;
sine[38717]=-56;
sine[38718]=-56;
sine[38719]=-56;
sine[38720]=-56;
sine[38721]=-56;
sine[38722]=-56;
sine[38723]=-56;
sine[38724]=-56;
sine[38725]=-56;
sine[38726]=-56;
sine[38727]=-56;
sine[38728]=-56;
sine[38729]=-56;
sine[38730]=-56;
sine[38731]=-56;
sine[38732]=-56;
sine[38733]=-56;
sine[38734]=-56;
sine[38735]=-56;
sine[38736]=-56;
sine[38737]=-56;
sine[38738]=-56;
sine[38739]=-56;
sine[38740]=-56;
sine[38741]=-56;
sine[38742]=-56;
sine[38743]=-55;
sine[38744]=-55;
sine[38745]=-55;
sine[38746]=-55;
sine[38747]=-55;
sine[38748]=-55;
sine[38749]=-55;
sine[38750]=-55;
sine[38751]=-55;
sine[38752]=-55;
sine[38753]=-55;
sine[38754]=-55;
sine[38755]=-55;
sine[38756]=-55;
sine[38757]=-55;
sine[38758]=-55;
sine[38759]=-55;
sine[38760]=-55;
sine[38761]=-55;
sine[38762]=-55;
sine[38763]=-55;
sine[38764]=-55;
sine[38765]=-55;
sine[38766]=-55;
sine[38767]=-55;
sine[38768]=-55;
sine[38769]=-55;
sine[38770]=-55;
sine[38771]=-55;
sine[38772]=-54;
sine[38773]=-54;
sine[38774]=-54;
sine[38775]=-54;
sine[38776]=-54;
sine[38777]=-54;
sine[38778]=-54;
sine[38779]=-54;
sine[38780]=-54;
sine[38781]=-54;
sine[38782]=-54;
sine[38783]=-54;
sine[38784]=-54;
sine[38785]=-54;
sine[38786]=-54;
sine[38787]=-54;
sine[38788]=-54;
sine[38789]=-54;
sine[38790]=-54;
sine[38791]=-54;
sine[38792]=-54;
sine[38793]=-54;
sine[38794]=-54;
sine[38795]=-54;
sine[38796]=-54;
sine[38797]=-54;
sine[38798]=-54;
sine[38799]=-54;
sine[38800]=-53;
sine[38801]=-53;
sine[38802]=-53;
sine[38803]=-53;
sine[38804]=-53;
sine[38805]=-53;
sine[38806]=-53;
sine[38807]=-53;
sine[38808]=-53;
sine[38809]=-53;
sine[38810]=-53;
sine[38811]=-53;
sine[38812]=-53;
sine[38813]=-53;
sine[38814]=-53;
sine[38815]=-53;
sine[38816]=-53;
sine[38817]=-53;
sine[38818]=-53;
sine[38819]=-53;
sine[38820]=-53;
sine[38821]=-53;
sine[38822]=-53;
sine[38823]=-53;
sine[38824]=-53;
sine[38825]=-53;
sine[38826]=-53;
sine[38827]=-53;
sine[38828]=-52;
sine[38829]=-52;
sine[38830]=-52;
sine[38831]=-52;
sine[38832]=-52;
sine[38833]=-52;
sine[38834]=-52;
sine[38835]=-52;
sine[38836]=-52;
sine[38837]=-52;
sine[38838]=-52;
sine[38839]=-52;
sine[38840]=-52;
sine[38841]=-52;
sine[38842]=-52;
sine[38843]=-52;
sine[38844]=-52;
sine[38845]=-52;
sine[38846]=-52;
sine[38847]=-52;
sine[38848]=-52;
sine[38849]=-52;
sine[38850]=-52;
sine[38851]=-52;
sine[38852]=-52;
sine[38853]=-52;
sine[38854]=-52;
sine[38855]=-51;
sine[38856]=-51;
sine[38857]=-51;
sine[38858]=-51;
sine[38859]=-51;
sine[38860]=-51;
sine[38861]=-51;
sine[38862]=-51;
sine[38863]=-51;
sine[38864]=-51;
sine[38865]=-51;
sine[38866]=-51;
sine[38867]=-51;
sine[38868]=-51;
sine[38869]=-51;
sine[38870]=-51;
sine[38871]=-51;
sine[38872]=-51;
sine[38873]=-51;
sine[38874]=-51;
sine[38875]=-51;
sine[38876]=-51;
sine[38877]=-51;
sine[38878]=-51;
sine[38879]=-51;
sine[38880]=-51;
sine[38881]=-51;
sine[38882]=-50;
sine[38883]=-50;
sine[38884]=-50;
sine[38885]=-50;
sine[38886]=-50;
sine[38887]=-50;
sine[38888]=-50;
sine[38889]=-50;
sine[38890]=-50;
sine[38891]=-50;
sine[38892]=-50;
sine[38893]=-50;
sine[38894]=-50;
sine[38895]=-50;
sine[38896]=-50;
sine[38897]=-50;
sine[38898]=-50;
sine[38899]=-50;
sine[38900]=-50;
sine[38901]=-50;
sine[38902]=-50;
sine[38903]=-50;
sine[38904]=-50;
sine[38905]=-50;
sine[38906]=-50;
sine[38907]=-50;
sine[38908]=-49;
sine[38909]=-49;
sine[38910]=-49;
sine[38911]=-49;
sine[38912]=-49;
sine[38913]=-49;
sine[38914]=-49;
sine[38915]=-49;
sine[38916]=-49;
sine[38917]=-49;
sine[38918]=-49;
sine[38919]=-49;
sine[38920]=-49;
sine[38921]=-49;
sine[38922]=-49;
sine[38923]=-49;
sine[38924]=-49;
sine[38925]=-49;
sine[38926]=-49;
sine[38927]=-49;
sine[38928]=-49;
sine[38929]=-49;
sine[38930]=-49;
sine[38931]=-49;
sine[38932]=-49;
sine[38933]=-49;
sine[38934]=-49;
sine[38935]=-48;
sine[38936]=-48;
sine[38937]=-48;
sine[38938]=-48;
sine[38939]=-48;
sine[38940]=-48;
sine[38941]=-48;
sine[38942]=-48;
sine[38943]=-48;
sine[38944]=-48;
sine[38945]=-48;
sine[38946]=-48;
sine[38947]=-48;
sine[38948]=-48;
sine[38949]=-48;
sine[38950]=-48;
sine[38951]=-48;
sine[38952]=-48;
sine[38953]=-48;
sine[38954]=-48;
sine[38955]=-48;
sine[38956]=-48;
sine[38957]=-48;
sine[38958]=-48;
sine[38959]=-48;
sine[38960]=-47;
sine[38961]=-47;
sine[38962]=-47;
sine[38963]=-47;
sine[38964]=-47;
sine[38965]=-47;
sine[38966]=-47;
sine[38967]=-47;
sine[38968]=-47;
sine[38969]=-47;
sine[38970]=-47;
sine[38971]=-47;
sine[38972]=-47;
sine[38973]=-47;
sine[38974]=-47;
sine[38975]=-47;
sine[38976]=-47;
sine[38977]=-47;
sine[38978]=-47;
sine[38979]=-47;
sine[38980]=-47;
sine[38981]=-47;
sine[38982]=-47;
sine[38983]=-47;
sine[38984]=-47;
sine[38985]=-47;
sine[38986]=-46;
sine[38987]=-46;
sine[38988]=-46;
sine[38989]=-46;
sine[38990]=-46;
sine[38991]=-46;
sine[38992]=-46;
sine[38993]=-46;
sine[38994]=-46;
sine[38995]=-46;
sine[38996]=-46;
sine[38997]=-46;
sine[38998]=-46;
sine[38999]=-46;
sine[39000]=-46;
sine[39001]=-46;
sine[39002]=-46;
sine[39003]=-46;
sine[39004]=-46;
sine[39005]=-46;
sine[39006]=-46;
sine[39007]=-46;
sine[39008]=-46;
sine[39009]=-46;
sine[39010]=-46;
sine[39011]=-45;
sine[39012]=-45;
sine[39013]=-45;
sine[39014]=-45;
sine[39015]=-45;
sine[39016]=-45;
sine[39017]=-45;
sine[39018]=-45;
sine[39019]=-45;
sine[39020]=-45;
sine[39021]=-45;
sine[39022]=-45;
sine[39023]=-45;
sine[39024]=-45;
sine[39025]=-45;
sine[39026]=-45;
sine[39027]=-45;
sine[39028]=-45;
sine[39029]=-45;
sine[39030]=-45;
sine[39031]=-45;
sine[39032]=-45;
sine[39033]=-45;
sine[39034]=-45;
sine[39035]=-45;
sine[39036]=-44;
sine[39037]=-44;
sine[39038]=-44;
sine[39039]=-44;
sine[39040]=-44;
sine[39041]=-44;
sine[39042]=-44;
sine[39043]=-44;
sine[39044]=-44;
sine[39045]=-44;
sine[39046]=-44;
sine[39047]=-44;
sine[39048]=-44;
sine[39049]=-44;
sine[39050]=-44;
sine[39051]=-44;
sine[39052]=-44;
sine[39053]=-44;
sine[39054]=-44;
sine[39055]=-44;
sine[39056]=-44;
sine[39057]=-44;
sine[39058]=-44;
sine[39059]=-44;
sine[39060]=-44;
sine[39061]=-43;
sine[39062]=-43;
sine[39063]=-43;
sine[39064]=-43;
sine[39065]=-43;
sine[39066]=-43;
sine[39067]=-43;
sine[39068]=-43;
sine[39069]=-43;
sine[39070]=-43;
sine[39071]=-43;
sine[39072]=-43;
sine[39073]=-43;
sine[39074]=-43;
sine[39075]=-43;
sine[39076]=-43;
sine[39077]=-43;
sine[39078]=-43;
sine[39079]=-43;
sine[39080]=-43;
sine[39081]=-43;
sine[39082]=-43;
sine[39083]=-43;
sine[39084]=-43;
sine[39085]=-42;
sine[39086]=-42;
sine[39087]=-42;
sine[39088]=-42;
sine[39089]=-42;
sine[39090]=-42;
sine[39091]=-42;
sine[39092]=-42;
sine[39093]=-42;
sine[39094]=-42;
sine[39095]=-42;
sine[39096]=-42;
sine[39097]=-42;
sine[39098]=-42;
sine[39099]=-42;
sine[39100]=-42;
sine[39101]=-42;
sine[39102]=-42;
sine[39103]=-42;
sine[39104]=-42;
sine[39105]=-42;
sine[39106]=-42;
sine[39107]=-42;
sine[39108]=-42;
sine[39109]=-41;
sine[39110]=-41;
sine[39111]=-41;
sine[39112]=-41;
sine[39113]=-41;
sine[39114]=-41;
sine[39115]=-41;
sine[39116]=-41;
sine[39117]=-41;
sine[39118]=-41;
sine[39119]=-41;
sine[39120]=-41;
sine[39121]=-41;
sine[39122]=-41;
sine[39123]=-41;
sine[39124]=-41;
sine[39125]=-41;
sine[39126]=-41;
sine[39127]=-41;
sine[39128]=-41;
sine[39129]=-41;
sine[39130]=-41;
sine[39131]=-41;
sine[39132]=-41;
sine[39133]=-40;
sine[39134]=-40;
sine[39135]=-40;
sine[39136]=-40;
sine[39137]=-40;
sine[39138]=-40;
sine[39139]=-40;
sine[39140]=-40;
sine[39141]=-40;
sine[39142]=-40;
sine[39143]=-40;
sine[39144]=-40;
sine[39145]=-40;
sine[39146]=-40;
sine[39147]=-40;
sine[39148]=-40;
sine[39149]=-40;
sine[39150]=-40;
sine[39151]=-40;
sine[39152]=-40;
sine[39153]=-40;
sine[39154]=-40;
sine[39155]=-40;
sine[39156]=-40;
sine[39157]=-39;
sine[39158]=-39;
sine[39159]=-39;
sine[39160]=-39;
sine[39161]=-39;
sine[39162]=-39;
sine[39163]=-39;
sine[39164]=-39;
sine[39165]=-39;
sine[39166]=-39;
sine[39167]=-39;
sine[39168]=-39;
sine[39169]=-39;
sine[39170]=-39;
sine[39171]=-39;
sine[39172]=-39;
sine[39173]=-39;
sine[39174]=-39;
sine[39175]=-39;
sine[39176]=-39;
sine[39177]=-39;
sine[39178]=-39;
sine[39179]=-39;
sine[39180]=-38;
sine[39181]=-38;
sine[39182]=-38;
sine[39183]=-38;
sine[39184]=-38;
sine[39185]=-38;
sine[39186]=-38;
sine[39187]=-38;
sine[39188]=-38;
sine[39189]=-38;
sine[39190]=-38;
sine[39191]=-38;
sine[39192]=-38;
sine[39193]=-38;
sine[39194]=-38;
sine[39195]=-38;
sine[39196]=-38;
sine[39197]=-38;
sine[39198]=-38;
sine[39199]=-38;
sine[39200]=-38;
sine[39201]=-38;
sine[39202]=-38;
sine[39203]=-38;
sine[39204]=-37;
sine[39205]=-37;
sine[39206]=-37;
sine[39207]=-37;
sine[39208]=-37;
sine[39209]=-37;
sine[39210]=-37;
sine[39211]=-37;
sine[39212]=-37;
sine[39213]=-37;
sine[39214]=-37;
sine[39215]=-37;
sine[39216]=-37;
sine[39217]=-37;
sine[39218]=-37;
sine[39219]=-37;
sine[39220]=-37;
sine[39221]=-37;
sine[39222]=-37;
sine[39223]=-37;
sine[39224]=-37;
sine[39225]=-37;
sine[39226]=-37;
sine[39227]=-36;
sine[39228]=-36;
sine[39229]=-36;
sine[39230]=-36;
sine[39231]=-36;
sine[39232]=-36;
sine[39233]=-36;
sine[39234]=-36;
sine[39235]=-36;
sine[39236]=-36;
sine[39237]=-36;
sine[39238]=-36;
sine[39239]=-36;
sine[39240]=-36;
sine[39241]=-36;
sine[39242]=-36;
sine[39243]=-36;
sine[39244]=-36;
sine[39245]=-36;
sine[39246]=-36;
sine[39247]=-36;
sine[39248]=-36;
sine[39249]=-36;
sine[39250]=-35;
sine[39251]=-35;
sine[39252]=-35;
sine[39253]=-35;
sine[39254]=-35;
sine[39255]=-35;
sine[39256]=-35;
sine[39257]=-35;
sine[39258]=-35;
sine[39259]=-35;
sine[39260]=-35;
sine[39261]=-35;
sine[39262]=-35;
sine[39263]=-35;
sine[39264]=-35;
sine[39265]=-35;
sine[39266]=-35;
sine[39267]=-35;
sine[39268]=-35;
sine[39269]=-35;
sine[39270]=-35;
sine[39271]=-35;
sine[39272]=-35;
sine[39273]=-34;
sine[39274]=-34;
sine[39275]=-34;
sine[39276]=-34;
sine[39277]=-34;
sine[39278]=-34;
sine[39279]=-34;
sine[39280]=-34;
sine[39281]=-34;
sine[39282]=-34;
sine[39283]=-34;
sine[39284]=-34;
sine[39285]=-34;
sine[39286]=-34;
sine[39287]=-34;
sine[39288]=-34;
sine[39289]=-34;
sine[39290]=-34;
sine[39291]=-34;
sine[39292]=-34;
sine[39293]=-34;
sine[39294]=-34;
sine[39295]=-33;
sine[39296]=-33;
sine[39297]=-33;
sine[39298]=-33;
sine[39299]=-33;
sine[39300]=-33;
sine[39301]=-33;
sine[39302]=-33;
sine[39303]=-33;
sine[39304]=-33;
sine[39305]=-33;
sine[39306]=-33;
sine[39307]=-33;
sine[39308]=-33;
sine[39309]=-33;
sine[39310]=-33;
sine[39311]=-33;
sine[39312]=-33;
sine[39313]=-33;
sine[39314]=-33;
sine[39315]=-33;
sine[39316]=-33;
sine[39317]=-33;
sine[39318]=-32;
sine[39319]=-32;
sine[39320]=-32;
sine[39321]=-32;
sine[39322]=-32;
sine[39323]=-32;
sine[39324]=-32;
sine[39325]=-32;
sine[39326]=-32;
sine[39327]=-32;
sine[39328]=-32;
sine[39329]=-32;
sine[39330]=-32;
sine[39331]=-32;
sine[39332]=-32;
sine[39333]=-32;
sine[39334]=-32;
sine[39335]=-32;
sine[39336]=-32;
sine[39337]=-32;
sine[39338]=-32;
sine[39339]=-32;
sine[39340]=-31;
sine[39341]=-31;
sine[39342]=-31;
sine[39343]=-31;
sine[39344]=-31;
sine[39345]=-31;
sine[39346]=-31;
sine[39347]=-31;
sine[39348]=-31;
sine[39349]=-31;
sine[39350]=-31;
sine[39351]=-31;
sine[39352]=-31;
sine[39353]=-31;
sine[39354]=-31;
sine[39355]=-31;
sine[39356]=-31;
sine[39357]=-31;
sine[39358]=-31;
sine[39359]=-31;
sine[39360]=-31;
sine[39361]=-31;
sine[39362]=-30;
sine[39363]=-30;
sine[39364]=-30;
sine[39365]=-30;
sine[39366]=-30;
sine[39367]=-30;
sine[39368]=-30;
sine[39369]=-30;
sine[39370]=-30;
sine[39371]=-30;
sine[39372]=-30;
sine[39373]=-30;
sine[39374]=-30;
sine[39375]=-30;
sine[39376]=-30;
sine[39377]=-30;
sine[39378]=-30;
sine[39379]=-30;
sine[39380]=-30;
sine[39381]=-30;
sine[39382]=-30;
sine[39383]=-30;
sine[39384]=-29;
sine[39385]=-29;
sine[39386]=-29;
sine[39387]=-29;
sine[39388]=-29;
sine[39389]=-29;
sine[39390]=-29;
sine[39391]=-29;
sine[39392]=-29;
sine[39393]=-29;
sine[39394]=-29;
sine[39395]=-29;
sine[39396]=-29;
sine[39397]=-29;
sine[39398]=-29;
sine[39399]=-29;
sine[39400]=-29;
sine[39401]=-29;
sine[39402]=-29;
sine[39403]=-29;
sine[39404]=-29;
sine[39405]=-29;
sine[39406]=-28;
sine[39407]=-28;
sine[39408]=-28;
sine[39409]=-28;
sine[39410]=-28;
sine[39411]=-28;
sine[39412]=-28;
sine[39413]=-28;
sine[39414]=-28;
sine[39415]=-28;
sine[39416]=-28;
sine[39417]=-28;
sine[39418]=-28;
sine[39419]=-28;
sine[39420]=-28;
sine[39421]=-28;
sine[39422]=-28;
sine[39423]=-28;
sine[39424]=-28;
sine[39425]=-28;
sine[39426]=-28;
sine[39427]=-28;
sine[39428]=-27;
sine[39429]=-27;
sine[39430]=-27;
sine[39431]=-27;
sine[39432]=-27;
sine[39433]=-27;
sine[39434]=-27;
sine[39435]=-27;
sine[39436]=-27;
sine[39437]=-27;
sine[39438]=-27;
sine[39439]=-27;
sine[39440]=-27;
sine[39441]=-27;
sine[39442]=-27;
sine[39443]=-27;
sine[39444]=-27;
sine[39445]=-27;
sine[39446]=-27;
sine[39447]=-27;
sine[39448]=-27;
sine[39449]=-27;
sine[39450]=-26;
sine[39451]=-26;
sine[39452]=-26;
sine[39453]=-26;
sine[39454]=-26;
sine[39455]=-26;
sine[39456]=-26;
sine[39457]=-26;
sine[39458]=-26;
sine[39459]=-26;
sine[39460]=-26;
sine[39461]=-26;
sine[39462]=-26;
sine[39463]=-26;
sine[39464]=-26;
sine[39465]=-26;
sine[39466]=-26;
sine[39467]=-26;
sine[39468]=-26;
sine[39469]=-26;
sine[39470]=-26;
sine[39471]=-25;
sine[39472]=-25;
sine[39473]=-25;
sine[39474]=-25;
sine[39475]=-25;
sine[39476]=-25;
sine[39477]=-25;
sine[39478]=-25;
sine[39479]=-25;
sine[39480]=-25;
sine[39481]=-25;
sine[39482]=-25;
sine[39483]=-25;
sine[39484]=-25;
sine[39485]=-25;
sine[39486]=-25;
sine[39487]=-25;
sine[39488]=-25;
sine[39489]=-25;
sine[39490]=-25;
sine[39491]=-25;
sine[39492]=-25;
sine[39493]=-24;
sine[39494]=-24;
sine[39495]=-24;
sine[39496]=-24;
sine[39497]=-24;
sine[39498]=-24;
sine[39499]=-24;
sine[39500]=-24;
sine[39501]=-24;
sine[39502]=-24;
sine[39503]=-24;
sine[39504]=-24;
sine[39505]=-24;
sine[39506]=-24;
sine[39507]=-24;
sine[39508]=-24;
sine[39509]=-24;
sine[39510]=-24;
sine[39511]=-24;
sine[39512]=-24;
sine[39513]=-24;
sine[39514]=-23;
sine[39515]=-23;
sine[39516]=-23;
sine[39517]=-23;
sine[39518]=-23;
sine[39519]=-23;
sine[39520]=-23;
sine[39521]=-23;
sine[39522]=-23;
sine[39523]=-23;
sine[39524]=-23;
sine[39525]=-23;
sine[39526]=-23;
sine[39527]=-23;
sine[39528]=-23;
sine[39529]=-23;
sine[39530]=-23;
sine[39531]=-23;
sine[39532]=-23;
sine[39533]=-23;
sine[39534]=-23;
sine[39535]=-23;
sine[39536]=-22;
sine[39537]=-22;
sine[39538]=-22;
sine[39539]=-22;
sine[39540]=-22;
sine[39541]=-22;
sine[39542]=-22;
sine[39543]=-22;
sine[39544]=-22;
sine[39545]=-22;
sine[39546]=-22;
sine[39547]=-22;
sine[39548]=-22;
sine[39549]=-22;
sine[39550]=-22;
sine[39551]=-22;
sine[39552]=-22;
sine[39553]=-22;
sine[39554]=-22;
sine[39555]=-22;
sine[39556]=-22;
sine[39557]=-21;
sine[39558]=-21;
sine[39559]=-21;
sine[39560]=-21;
sine[39561]=-21;
sine[39562]=-21;
sine[39563]=-21;
sine[39564]=-21;
sine[39565]=-21;
sine[39566]=-21;
sine[39567]=-21;
sine[39568]=-21;
sine[39569]=-21;
sine[39570]=-21;
sine[39571]=-21;
sine[39572]=-21;
sine[39573]=-21;
sine[39574]=-21;
sine[39575]=-21;
sine[39576]=-21;
sine[39577]=-21;
sine[39578]=-20;
sine[39579]=-20;
sine[39580]=-20;
sine[39581]=-20;
sine[39582]=-20;
sine[39583]=-20;
sine[39584]=-20;
sine[39585]=-20;
sine[39586]=-20;
sine[39587]=-20;
sine[39588]=-20;
sine[39589]=-20;
sine[39590]=-20;
sine[39591]=-20;
sine[39592]=-20;
sine[39593]=-20;
sine[39594]=-20;
sine[39595]=-20;
sine[39596]=-20;
sine[39597]=-20;
sine[39598]=-20;
sine[39599]=-19;
sine[39600]=-19;
sine[39601]=-19;
sine[39602]=-19;
sine[39603]=-19;
sine[39604]=-19;
sine[39605]=-19;
sine[39606]=-19;
sine[39607]=-19;
sine[39608]=-19;
sine[39609]=-19;
sine[39610]=-19;
sine[39611]=-19;
sine[39612]=-19;
sine[39613]=-19;
sine[39614]=-19;
sine[39615]=-19;
sine[39616]=-19;
sine[39617]=-19;
sine[39618]=-19;
sine[39619]=-19;
sine[39620]=-18;
sine[39621]=-18;
sine[39622]=-18;
sine[39623]=-18;
sine[39624]=-18;
sine[39625]=-18;
sine[39626]=-18;
sine[39627]=-18;
sine[39628]=-18;
sine[39629]=-18;
sine[39630]=-18;
sine[39631]=-18;
sine[39632]=-18;
sine[39633]=-18;
sine[39634]=-18;
sine[39635]=-18;
sine[39636]=-18;
sine[39637]=-18;
sine[39638]=-18;
sine[39639]=-18;
sine[39640]=-18;
sine[39641]=-17;
sine[39642]=-17;
sine[39643]=-17;
sine[39644]=-17;
sine[39645]=-17;
sine[39646]=-17;
sine[39647]=-17;
sine[39648]=-17;
sine[39649]=-17;
sine[39650]=-17;
sine[39651]=-17;
sine[39652]=-17;
sine[39653]=-17;
sine[39654]=-17;
sine[39655]=-17;
sine[39656]=-17;
sine[39657]=-17;
sine[39658]=-17;
sine[39659]=-17;
sine[39660]=-17;
sine[39661]=-17;
sine[39662]=-16;
sine[39663]=-16;
sine[39664]=-16;
sine[39665]=-16;
sine[39666]=-16;
sine[39667]=-16;
sine[39668]=-16;
sine[39669]=-16;
sine[39670]=-16;
sine[39671]=-16;
sine[39672]=-16;
sine[39673]=-16;
sine[39674]=-16;
sine[39675]=-16;
sine[39676]=-16;
sine[39677]=-16;
sine[39678]=-16;
sine[39679]=-16;
sine[39680]=-16;
sine[39681]=-16;
sine[39682]=-16;
sine[39683]=-15;
sine[39684]=-15;
sine[39685]=-15;
sine[39686]=-15;
sine[39687]=-15;
sine[39688]=-15;
sine[39689]=-15;
sine[39690]=-15;
sine[39691]=-15;
sine[39692]=-15;
sine[39693]=-15;
sine[39694]=-15;
sine[39695]=-15;
sine[39696]=-15;
sine[39697]=-15;
sine[39698]=-15;
sine[39699]=-15;
sine[39700]=-15;
sine[39701]=-15;
sine[39702]=-15;
sine[39703]=-14;
sine[39704]=-14;
sine[39705]=-14;
sine[39706]=-14;
sine[39707]=-14;
sine[39708]=-14;
sine[39709]=-14;
sine[39710]=-14;
sine[39711]=-14;
sine[39712]=-14;
sine[39713]=-14;
sine[39714]=-14;
sine[39715]=-14;
sine[39716]=-14;
sine[39717]=-14;
sine[39718]=-14;
sine[39719]=-14;
sine[39720]=-14;
sine[39721]=-14;
sine[39722]=-14;
sine[39723]=-14;
sine[39724]=-13;
sine[39725]=-13;
sine[39726]=-13;
sine[39727]=-13;
sine[39728]=-13;
sine[39729]=-13;
sine[39730]=-13;
sine[39731]=-13;
sine[39732]=-13;
sine[39733]=-13;
sine[39734]=-13;
sine[39735]=-13;
sine[39736]=-13;
sine[39737]=-13;
sine[39738]=-13;
sine[39739]=-13;
sine[39740]=-13;
sine[39741]=-13;
sine[39742]=-13;
sine[39743]=-13;
sine[39744]=-13;
sine[39745]=-12;
sine[39746]=-12;
sine[39747]=-12;
sine[39748]=-12;
sine[39749]=-12;
sine[39750]=-12;
sine[39751]=-12;
sine[39752]=-12;
sine[39753]=-12;
sine[39754]=-12;
sine[39755]=-12;
sine[39756]=-12;
sine[39757]=-12;
sine[39758]=-12;
sine[39759]=-12;
sine[39760]=-12;
sine[39761]=-12;
sine[39762]=-12;
sine[39763]=-12;
sine[39764]=-12;
sine[39765]=-11;
sine[39766]=-11;
sine[39767]=-11;
sine[39768]=-11;
sine[39769]=-11;
sine[39770]=-11;
sine[39771]=-11;
sine[39772]=-11;
sine[39773]=-11;
sine[39774]=-11;
sine[39775]=-11;
sine[39776]=-11;
sine[39777]=-11;
sine[39778]=-11;
sine[39779]=-11;
sine[39780]=-11;
sine[39781]=-11;
sine[39782]=-11;
sine[39783]=-11;
sine[39784]=-11;
sine[39785]=-11;
sine[39786]=-10;
sine[39787]=-10;
sine[39788]=-10;
sine[39789]=-10;
sine[39790]=-10;
sine[39791]=-10;
sine[39792]=-10;
sine[39793]=-10;
sine[39794]=-10;
sine[39795]=-10;
sine[39796]=-10;
sine[39797]=-10;
sine[39798]=-10;
sine[39799]=-10;
sine[39800]=-10;
sine[39801]=-10;
sine[39802]=-10;
sine[39803]=-10;
sine[39804]=-10;
sine[39805]=-10;
sine[39806]=-9;
sine[39807]=-9;
sine[39808]=-9;
sine[39809]=-9;
sine[39810]=-9;
sine[39811]=-9;
sine[39812]=-9;
sine[39813]=-9;
sine[39814]=-9;
sine[39815]=-9;
sine[39816]=-9;
sine[39817]=-9;
sine[39818]=-9;
sine[39819]=-9;
sine[39820]=-9;
sine[39821]=-9;
sine[39822]=-9;
sine[39823]=-9;
sine[39824]=-9;
sine[39825]=-9;
sine[39826]=-9;
sine[39827]=-8;
sine[39828]=-8;
sine[39829]=-8;
sine[39830]=-8;
sine[39831]=-8;
sine[39832]=-8;
sine[39833]=-8;
sine[39834]=-8;
sine[39835]=-8;
sine[39836]=-8;
sine[39837]=-8;
sine[39838]=-8;
sine[39839]=-8;
sine[39840]=-8;
sine[39841]=-8;
sine[39842]=-8;
sine[39843]=-8;
sine[39844]=-8;
sine[39845]=-8;
sine[39846]=-8;
sine[39847]=-7;
sine[39848]=-7;
sine[39849]=-7;
sine[39850]=-7;
sine[39851]=-7;
sine[39852]=-7;
sine[39853]=-7;
sine[39854]=-7;
sine[39855]=-7;
sine[39856]=-7;
sine[39857]=-7;
sine[39858]=-7;
sine[39859]=-7;
sine[39860]=-7;
sine[39861]=-7;
sine[39862]=-7;
sine[39863]=-7;
sine[39864]=-7;
sine[39865]=-7;
sine[39866]=-7;
sine[39867]=-7;
sine[39868]=-6;
sine[39869]=-6;
sine[39870]=-6;
sine[39871]=-6;
sine[39872]=-6;
sine[39873]=-6;
sine[39874]=-6;
sine[39875]=-6;
sine[39876]=-6;
sine[39877]=-6;
sine[39878]=-6;
sine[39879]=-6;
sine[39880]=-6;
sine[39881]=-6;
sine[39882]=-6;
sine[39883]=-6;
sine[39884]=-6;
sine[39885]=-6;
sine[39886]=-6;
sine[39887]=-6;
sine[39888]=-5;
sine[39889]=-5;
sine[39890]=-5;
sine[39891]=-5;
sine[39892]=-5;
sine[39893]=-5;
sine[39894]=-5;
sine[39895]=-5;
sine[39896]=-5;
sine[39897]=-5;
sine[39898]=-5;
sine[39899]=-5;
sine[39900]=-5;
sine[39901]=-5;
sine[39902]=-5;
sine[39903]=-5;
sine[39904]=-5;
sine[39905]=-5;
sine[39906]=-5;
sine[39907]=-5;
sine[39908]=-5;
sine[39909]=-4;
sine[39910]=-4;
sine[39911]=-4;
sine[39912]=-4;
sine[39913]=-4;
sine[39914]=-4;
sine[39915]=-4;
sine[39916]=-4;
sine[39917]=-4;
sine[39918]=-4;
sine[39919]=-4;
sine[39920]=-4;
sine[39921]=-4;
sine[39922]=-4;
sine[39923]=-4;
sine[39924]=-4;
sine[39925]=-4;
sine[39926]=-4;
sine[39927]=-4;
sine[39928]=-4;
sine[39929]=-3;
sine[39930]=-3;
sine[39931]=-3;
sine[39932]=-3;
sine[39933]=-3;
sine[39934]=-3;
sine[39935]=-3;
sine[39936]=-3;
sine[39937]=-3;
sine[39938]=-3;
sine[39939]=-3;
sine[39940]=-3;
sine[39941]=-3;
sine[39942]=-3;
sine[39943]=-3;
sine[39944]=-3;
sine[39945]=-3;
sine[39946]=-3;
sine[39947]=-3;
sine[39948]=-3;
sine[39949]=-3;
sine[39950]=-2;
sine[39951]=-2;
sine[39952]=-2;
sine[39953]=-2;
sine[39954]=-2;
sine[39955]=-2;
sine[39956]=-2;
sine[39957]=-2;
sine[39958]=-2;
sine[39959]=-2;
sine[39960]=-2;
sine[39961]=-2;
sine[39962]=-2;
sine[39963]=-2;
sine[39964]=-2;
sine[39965]=-2;
sine[39966]=-2;
sine[39967]=-2;
sine[39968]=-2;
sine[39969]=-2;
sine[39970]=-1;
sine[39971]=-1;
sine[39972]=-1;
sine[39973]=-1;
sine[39974]=-1;
sine[39975]=-1;
sine[39976]=-1;
sine[39977]=-1;
sine[39978]=-1;
sine[39979]=-1;
sine[39980]=-1;
sine[39981]=-1;
sine[39982]=-1;
sine[39983]=-1;
sine[39984]=-1;
sine[39985]=-1;
sine[39986]=-1;
sine[39987]=-1;
sine[39988]=-1;
sine[39989]=-1;
sine[39990]=0;
sine[39991]=0;
sine[39992]=0;
sine[39993]=0;
sine[39994]=0;
sine[39995]=0;
sine[39996]=0;
sine[39997]=0;
sine[39998]=0;
sine[39999]=0;
sine[40000]=0;




    end
    
    
    always@ (posedge(Clk))
    begin
        sine_out = sine[i];
        cos_out=cos[i];
        i = i+ 1;
        if(i == 40000)
            i = 0;
    end

endmodule
